module AsyncFifo(input ulpi_clk, input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [7:0] io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output[7:0] io_deq_bits
    //output[4:0] io_count
);

  wire[7:0] T1;
  reg [7:0] mem [15:0];
  wire[7:0] T2;
  wire T3;
  wire[3:0] T4;
  reg [4:0] wptr_bin;
  wire[4:0] T20;
  wire[4:0] wptr_bin_next;
  wire[4:0] T21;
  wire T5;
  reg  not_full;
  wire T22;
  wire T6;
  wire T7;
  reg  s2_rst_deq;
  wire T23;
  reg  s1_rst_deq;
  wire T24;
  wire not_full_next;
  wire T8;
  wire[4:0] T9;
  wire[2:0] T10;
  reg [4:0] s2_rptr_gray;
  wire[4:0] T25;
  reg [4:0] s1_rptr_gray;
  wire[4:0] T26;
  reg [4:0] rptr_gray;
  wire[4:0] T27;
  wire[4:0] rptr_gray_next;
  wire[4:0] rptr_bin_next;
  wire[4:0] T28;
  wire T11;
  reg  not_empty;
  wire T29;
  wire T12;
  wire T13;
  reg  s2_rst_enq;
  wire T30;
  reg  s1_rst_enq;
  wire T31;
  wire not_empty_next;
  wire T14;
  reg [4:0] s2_wptr_gray;
  wire[4:0] T32;
  reg [4:0] s1_wptr_gray;
  wire[4:0] T33;
  reg [4:0] wptr_gray;
  wire[4:0] T34;
  reg [4:0] rptr_bin;
  wire[4:0] T35;
  wire[4:0] T36;
  wire[3:0] T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire[4:0] wptr_gray_next;
  wire[4:0] T37;
  wire[3:0] T18;
  wire[3:0] T19;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 16; initvar = initvar+1)
      mem[initvar] = {1{$random}};
    wptr_bin = {1{$random}};
    not_full = {1{$random}};
    s2_rst_deq = {1{$random}};
    s1_rst_deq = {1{$random}};
    s2_rptr_gray = {1{$random}};
    s1_rptr_gray = {1{$random}};
    rptr_gray = {1{$random}};
    not_empty = {1{$random}};
    s2_rst_enq = {1{$random}};
    s1_rst_enq = {1{$random}};
    s2_wptr_gray = {1{$random}};
    s1_wptr_gray = {1{$random}};
    wptr_gray = {1{$random}};
    rptr_bin = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_count = {1{$random}};
// synthesis translate_on
`endif
  assign io_deq_bits = T1;
  assign T1 = mem[T19];
  assign T3 = io_enq_valid & io_enq_ready;
  assign T4 = wptr_bin[3:0];
  assign T20 = reset ? 5'h0 : wptr_bin_next;
  assign wptr_bin_next = wptr_bin + T21;
  assign T21 = {4'h0, T5};
  assign T5 = io_enq_valid & not_full;
  assign T22 = reset ? 1'h0 : T6;
  assign T6 = not_full_next & T7;
  assign T7 = s2_rst_deq ^ 1'h1;
  assign T23 = reset ? 1'h0 : s1_rst_deq;
  assign T24 = reset ? 1'h0 : reset;
  assign not_full_next = T8 ^ 1'h1;
  assign T8 = wptr_gray_next == T9;
  assign T9 = {T16, T10};
  assign T10 = s2_rptr_gray[2:0];
  assign T25 = reset ? 5'h0 : s1_rptr_gray;
  assign T26 = reset ? 5'h0 : rptr_gray;
  assign T27 = reset ? 5'h0 : rptr_gray_next;
  assign rptr_gray_next = T36 ^ rptr_bin_next;
  assign rptr_bin_next = rptr_bin + T28;
  assign T28 = {4'h0, T11};
  assign T11 = io_deq_ready & not_empty;
  assign T29 = reset ? 1'h0 : T12;
  assign T12 = not_empty_next & T13;
  assign T13 = s2_rst_enq ^ 1'h1;
  assign T30 = reset ? 1'h0 : s1_rst_enq;
  assign T31 = reset ? 1'h0 : reset;
  assign not_empty_next = T14 ^ 1'h1;
  assign T14 = rptr_gray_next == s2_wptr_gray;
  assign T32 = reset ? 5'h0 : s1_wptr_gray;
  assign T33 = reset ? 5'h0 : wptr_gray;
  assign T34 = reset ? 5'h0 : wptr_gray_next;
  assign T35 = reset ? 5'h0 : rptr_bin_next;
  assign T36 = {1'h0, T15};
  assign T15 = rptr_bin_next >> 1'h1;
  assign T16 = ~ T17;
  assign T17 = s2_rptr_gray[4:3];
  assign wptr_gray_next = T37 ^ wptr_bin_next;
  assign T37 = {1'h0, T18};
  assign T18 = wptr_bin_next >> 1'h1;
  assign T19 = rptr_bin[3:0];
  assign io_deq_valid = not_empty;
  assign io_enq_ready = not_full;

  always @(posedge ulpi_clk) begin
    if (T3)
      mem[T4] <= io_enq_bits;
    if(reset) begin
      wptr_bin <= 5'h0;
    end else begin
      wptr_bin <= wptr_bin_next;
    end
    if(reset) begin
      not_full <= 1'h0;
    end else begin
      not_full <= T6;
    end
    if(reset) begin
      s2_rst_deq <= 1'h0;
    end else begin
      s2_rst_deq <= s1_rst_deq;
    end
    if(reset) begin
      s1_rst_deq <= 1'h0;
    end else begin
      s1_rst_deq <= reset;
    end
    if(reset) begin
      s2_rptr_gray <= 5'h0;
    end else begin
      s2_rptr_gray <= s1_rptr_gray;
    end
    if(reset) begin
      s1_rptr_gray <= 5'h0;
    end else begin
      s1_rptr_gray <= rptr_gray;
    end
    if(reset) begin
      wptr_gray <= 5'h0;
    end else begin
      wptr_gray <= wptr_gray_next;
    end
  end
  always @(posedge clk) begin
    if(reset) begin
      rptr_gray <= 5'h0;
    end else begin
      rptr_gray <= rptr_gray_next;
    end
    if(reset) begin
      not_empty <= 1'h0;
    end else begin
      not_empty <= T12;
    end
    if(reset) begin
      s2_rst_enq <= 1'h0;
    end else begin
      s2_rst_enq <= s1_rst_enq;
    end
    if(reset) begin
      s1_rst_enq <= 1'h0;
    end else begin
      s1_rst_enq <= reset;
    end
    if(reset) begin
      s2_wptr_gray <= 5'h0;
    end else begin
      s2_wptr_gray <= s1_wptr_gray;
    end
    if(reset) begin
      s1_wptr_gray <= 5'h0;
    end else begin
      s1_wptr_gray <= wptr_gray;
    end
    if(reset) begin
      rptr_bin <= 5'h0;
    end else begin
      rptr_bin <= rptr_bin_next;
    end
  end
endmodule

module CounterWithNonBlockingReset(input clk, input reset,
    input  io_enable,
    input  io_rst,
    output[1:0] io_value
);

  reg [1:0] reg_;
  wire[1:0] T4;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] base;
  wire T3;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    reg_ = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = reg_;
  assign T4 = reset ? 2'h0 : T0;
  assign T0 = T3 ? reg_ : T1;
  assign T1 = io_enable ? T2 : reg_;
  assign T2 = base + 2'h1;
  assign base = io_rst ? 2'h0 : reg_;
  assign T3 = io_enable ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      reg_ <= 2'h0;
    end else if(T3) begin
      reg_ <= reg_;
    end else if(io_enable) begin
      reg_ <= T2;
    end
  end
endmodule

module WidthConverter(input clk, input reset,
    output io_wordIn_ready,
    input  io_wordIn_valid,
    input [7:0] io_wordIn_bits,
    input  io_wordOut_ready,
    output io_wordOut_valid,
    output[15:0] io_wordOut_bits
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire[15:0] T5;
  reg [7:0] R6;
  wire[7:0] T7;
  wire[7:0] T8;
  wire T9;
  reg [7:0] R10;
  wire[7:0] T11;
  wire[7:0] T12;
  wire[1:0] CounterWithNonBlockingReset_io_value;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R6 = {1{$random}};
    R10 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = T1 & io_wordOut_ready;
  assign T1 = CounterWithNonBlockingReset_io_value == 2'h2;
  assign T2 = T3 & io_wordIn_valid;
  assign T3 = T4 | io_wordOut_ready;
  assign T4 = T1 ^ 1'h1;
  assign io_wordOut_bits = T5;
  assign T5 = {R10, R6};
  assign T7 = T9 ? R6 : T8;
  assign T8 = T2 ? R10 : R6;
  assign T9 = T2 ^ 1'h1;
  assign T11 = T9 ? R10 : T12;
  assign T12 = T2 ? io_wordIn_bits : R10;
  assign io_wordOut_valid = T1;
  assign io_wordIn_ready = T3;
  CounterWithNonBlockingReset CounterWithNonBlockingReset(.clk(clk), .reset(reset),
       .io_enable( T2 ),
       .io_rst( T0 ),
       .io_value( CounterWithNonBlockingReset_io_value )
  );

  always @(posedge clk) begin
    if(T9) begin
      R6 <= R6;
    end else if(T2) begin
      R6 <= R10;
    end
    if(T9) begin
      R10 <= R10;
    end else if(T2) begin
      R10 <= io_wordIn_bits;
    end
  end
endmodule

module AsyncCounter_0(input clk, input reset,
    input  io_enable,
    output[7:0] io_value
);

  wire[7:0] T0;
  reg [7:0] v;
  wire[7:0] T5;
  wire[7:0] T1;
  wire[7:0] T2;
  wire[7:0] T3;
  wire T4;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    v = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = T0;
  assign T0 = io_enable ? T2 : v;
  assign T5 = reset ? 8'h0 : T1;
  assign T1 = io_enable ? T2 : v;
  assign T2 = T4 ? 8'h0 : T3;
  assign T3 = v + 8'h31;
  assign T4 = v == 8'h62;

  always @(posedge clk) begin
    if(reset) begin
      v <= 8'h0;
    end else if(io_enable) begin
      v <= T2;
    end
  end
endmodule

module CounterWithSyncAndAsyncReset_0(input clk, input reset,
    input  io_enable,
    input  io_syncRst,
    input  io_asyncRst,
    output[5:0] io_value
);

  wire[5:0] T0;
  reg [5:0] v;
  wire[5:0] T13;
  wire[5:0] T1;
  wire[5:0] T2;
  wire[5:0] T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire[5:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire[5:0] T12;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    v = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = T0;
  assign T0 = io_enable ? T12 : v;
  assign T13 = reset ? 6'h0 : T1;
  assign T1 = T9 ? T8 : T2;
  assign T2 = T5 ? 6'h0 : T3;
  assign T3 = T4 ? 6'h1 : v;
  assign T4 = io_enable & io_asyncRst;
  assign T5 = io_enable & T6;
  assign T6 = T7 & io_syncRst;
  assign T7 = io_asyncRst ^ 1'h1;
  assign T8 = v + 6'h1;
  assign T9 = io_enable & T10;
  assign T10 = T11 ^ 1'h1;
  assign T11 = io_asyncRst | io_syncRst;
  assign T12 = io_asyncRst ? 6'h0 : v;

  always @(posedge clk) begin
    if(reset) begin
      v <= 6'h0;
    end else if(T9) begin
      v <= T8;
    end else if(T5) begin
      v <= 6'h0;
    end else if(T4) begin
      v <= 6'h1;
    end
  end
endmodule

module CircularPeekQueue_0(input clk, input reset,
    input  io_writeEnable,
    input  io_nextBlock,
    input [15:0] io_input,
    output[15:0] io_output
);

  reg [7:0] writeAddr;
  wire[7:0] T10;
  wire[7:0] T0;
  wire[7:0] T1;
  wire T2;
  wire T3;
  wire[7:0] T4;
  wire T5;
  wire T6;
  wire[7:0] T7;
  wire[7:0] T11;
  wire[5:0] T8;
  wire T9;
  wire[7:0] currentBlockOffset_io_value;
  wire[5:0] inBlockReadOffset_io_value;
  wire[15:0] queue_b_dout;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    writeAddr = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T10 = reset ? 8'h31 : T0;
  assign T0 = T5 ? T4 : T1;
  assign T1 = T2 ? 8'h0 : writeAddr;
  assign T2 = io_writeEnable & T3;
  assign T3 = writeAddr == 8'h92;
  assign T4 = writeAddr + 8'h1;
  assign T5 = io_writeEnable & T6;
  assign T6 = T3 ^ 1'h1;
  assign T7 = currentBlockOffset_io_value + T11;
  assign T11 = {2'h0, T8};
  assign T8 = io_nextBlock ? 6'h0 : inBlockReadOffset_io_value;
  assign T9 = inBlockReadOffset_io_value == 6'h30;
  assign io_output = queue_b_dout;
  AsyncCounter_0 currentBlockOffset(.clk(clk), .reset(reset),
       .io_enable( io_nextBlock ),
       .io_value( currentBlockOffset_io_value )
  );
  CounterWithSyncAndAsyncReset_0 inBlockReadOffset(.clk(clk), .reset(reset),
       .io_enable( 1'h1 ),
       .io_syncRst( T9 ),
       .io_asyncRst( io_nextBlock ),
       .io_value( inBlockReadOffset_io_value )
  );
  DualPortBRAM # (
    .DATA(16),
    .ADDR(8)
  ) queue(.clk(clk),
       .b_addr( T7 ),
       //.b_din(  )
       .b_wr( 1'h0 ),
       .b_dout( queue_b_dout ),
       .a_addr( writeAddr ),
       .a_din( io_input ),
       .a_wr( io_writeEnable )
       //.a_dout(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign queue.b_din = {1{$random}};
// synthesis translate_on
`endif

  always @(posedge clk) begin
    if(reset) begin
      writeAddr <= 8'h31;
    end else if(T5) begin
      writeAddr <= T4;
    end else if(T2) begin
      writeAddr <= 8'h0;
    end
  end
endmodule

module Counter_0(input clk, input reset,
    input  io_enable,
    input  io_rst,
    output[5:0] io_value
);

  reg [5:0] v;
  wire[5:0] T6;
  wire[5:0] T0;
  wire[5:0] T1;
  wire T2;
  wire[5:0] T3;
  wire T4;
  wire T5;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    v = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = v;
  assign T6 = reset ? 6'h0 : T0;
  assign T0 = T4 ? T3 : T1;
  assign T1 = T2 ? 6'h0 : v;
  assign T2 = io_enable & io_rst;
  assign T3 = v + 6'h1;
  assign T4 = io_enable & T5;
  assign T5 = io_rst ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      v <= 6'h0;
    end else if(T4) begin
      v <= T3;
    end else if(T2) begin
      v <= 6'h0;
    end
  end
endmodule

module Counter_1(input clk, input reset,
    input  io_enable,
    input  io_rst,
    output[1:0] io_value
);

  reg [1:0] v;
  wire[1:0] T6;
  wire[1:0] T0;
  wire[1:0] T1;
  wire T2;
  wire[1:0] T3;
  wire T4;
  wire T5;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    v = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = v;
  assign T6 = reset ? 2'h0 : T0;
  assign T0 = T4 ? T3 : T1;
  assign T1 = T2 ? 2'h0 : v;
  assign T2 = io_enable & io_rst;
  assign T3 = v + 2'h1;
  assign T4 = io_enable & T5;
  assign T5 = io_rst ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      v <= 2'h0;
    end else if(T4) begin
      v <= T3;
    end else if(T2) begin
      v <= 2'h0;
    end
  end
endmodule

module UpDownCounter_0(input clk, input reset,
    input  io_up,
    input  io_down,
    output[1:0] io_value
);

  reg [1:0] reg_;
  wire[1:0] T10;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire T3;
  wire T4;
  wire T5;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    reg_ = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = reg_;
  assign T10 = reset ? 2'h0 : T0;
  assign T0 = T7 ? T6 : T1;
  assign T1 = T3 ? T2 : reg_;
  assign T2 = reg_ + 2'h1;
  assign T3 = T4 & io_up;
  assign T4 = T5 ^ 1'h1;
  assign T5 = io_up & io_down;
  assign T6 = reg_ - 2'h1;
  assign T7 = T8 & io_down;
  assign T8 = T9 ^ 1'h1;
  assign T9 = T5 | io_up;

  always @(posedge clk) begin
    if(reset) begin
      reg_ <= 2'h0;
    end else if(T7) begin
      reg_ <= T6;
    end else if(T3) begin
      reg_ <= T2;
    end
  end
endmodule

module Interleaver(input clk, input reset,
    output io_wordIn_ready,
    input  io_wordIn_valid,
    input [15:0] io_wordIn_bits,
    output[15:0] io_interleavedOut_3,
    output[15:0] io_interleavedOut_2,
    output[15:0] io_interleavedOut_1,
    output[15:0] io_interleavedOut_0,
    output io_startOut,
    input  io_pipeReady
);

  wire signalNewPeekBlock;
  wire T0;
  wire signalWritingLastWordInLastQueue;
  wire isLastQueue;
  wire signalWritingLastWord;
  wire isLastInputWordInBlock;
  wire signalReadingInput;
  wire isReady;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  reg  R9;
  wire T10;
  wire[5:0] wordCounter_io_value;
  wire[1:0] queueCounter_io_value;
  wire[1:0] readyBlocks_io_value;
  wire[15:0] CircularPeekQueue_io_output;
  wire[15:0] CircularPeekQueue_1_io_output;
  wire[15:0] CircularPeekQueue_2_io_output;
  wire[15:0] CircularPeekQueue_3_io_output;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R9 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign signalNewPeekBlock = io_pipeReady & T0;
  assign T0 = readyBlocks_io_value != 2'h0;
  assign signalWritingLastWordInLastQueue = signalWritingLastWord & isLastQueue;
  assign isLastQueue = queueCounter_io_value == 2'h3;
  assign signalWritingLastWord = signalReadingInput & isLastInputWordInBlock;
  assign isLastInputWordInBlock = wordCounter_io_value == 6'h30;
  assign signalReadingInput = io_wordIn_valid & isReady;
  assign isReady = readyBlocks_io_value != 2'h2;
  assign T1 = T2 & signalReadingInput;
  assign T2 = queueCounter_io_value == 2'h3;
  assign T3 = T4 & signalReadingInput;
  assign T4 = queueCounter_io_value == 2'h2;
  assign T5 = T6 & signalReadingInput;
  assign T6 = queueCounter_io_value == 2'h1;
  assign T7 = T8 & signalReadingInput;
  assign T8 = queueCounter_io_value == 2'h0;
  assign io_startOut = R9;
  assign T10 = reset ? 1'h0 : signalNewPeekBlock;
  assign io_interleavedOut_0 = CircularPeekQueue_io_output;
  assign io_interleavedOut_1 = CircularPeekQueue_1_io_output;
  assign io_interleavedOut_2 = CircularPeekQueue_2_io_output;
  assign io_interleavedOut_3 = CircularPeekQueue_3_io_output;
  assign io_wordIn_ready = isReady;
  CircularPeekQueue_0 CircularPeekQueue(.clk(clk), .reset(reset),
       .io_writeEnable( T7 ),
       .io_nextBlock( signalNewPeekBlock ),
       .io_input( io_wordIn_bits ),
       .io_output( CircularPeekQueue_io_output )
  );
  CircularPeekQueue_0 CircularPeekQueue_1(.clk(clk), .reset(reset),
       .io_writeEnable( T5 ),
       .io_nextBlock( signalNewPeekBlock ),
       .io_input( io_wordIn_bits ),
       .io_output( CircularPeekQueue_1_io_output )
  );
  CircularPeekQueue_0 CircularPeekQueue_2(.clk(clk), .reset(reset),
       .io_writeEnable( T3 ),
       .io_nextBlock( signalNewPeekBlock ),
       .io_input( io_wordIn_bits ),
       .io_output( CircularPeekQueue_2_io_output )
  );
  CircularPeekQueue_0 CircularPeekQueue_3(.clk(clk), .reset(reset),
       .io_writeEnable( T1 ),
       .io_nextBlock( signalNewPeekBlock ),
       .io_input( io_wordIn_bits ),
       .io_output( CircularPeekQueue_3_io_output )
  );
  Counter_0 wordCounter(.clk(clk), .reset(reset),
       .io_enable( signalReadingInput ),
       .io_rst( isLastInputWordInBlock ),
       .io_value( wordCounter_io_value )
  );
  Counter_1 queueCounter(.clk(clk), .reset(reset),
       .io_enable( signalWritingLastWord ),
       .io_rst( isLastQueue ),
       .io_value( queueCounter_io_value )
  );
  UpDownCounter_0 readyBlocks(.clk(clk), .reset(reset),
       .io_up( signalWritingLastWordInLastQueue ),
       .io_down( signalNewPeekBlock ),
       .io_value( readyBlocks_io_value )
  );

  always @(posedge clk) begin
    if(reset) begin
      R9 <= 1'h0;
    end else begin
      R9 <= signalNewPeekBlock;
    end
  end
endmodule

module Counter_3(input clk, input reset,
    input  io_enable,
    input  io_rst,
    output[8:0] io_value
);

  reg [8:0] v;
  wire[8:0] T6;
  wire[8:0] T0;
  wire[8:0] T1;
  wire T2;
  wire[8:0] T3;
  wire T4;
  wire T5;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    v = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = v;
  assign T6 = reset ? 9'h0 : T0;
  assign T0 = T4 ? T3 : T1;
  assign T1 = T2 ? 9'h0 : v;
  assign T2 = io_enable & io_rst;
  assign T3 = v + 9'h1;
  assign T4 = io_enable & T5;
  assign T5 = io_rst ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      v <= 9'h0;
    end else if(T4) begin
      v <= T3;
    end else if(T2) begin
      v <= 9'h0;
    end
  end
endmodule

module Counter_4(input clk, input reset,
    input  io_enable,
    input  io_rst,
    output[4:0] io_value
);

  reg [4:0] v;
  wire[4:0] T6;
  wire[4:0] T0;
  wire[4:0] T1;
  wire T2;
  wire[4:0] T3;
  wire T4;
  wire T5;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    v = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = v;
  assign T6 = reset ? 5'h0 : T0;
  assign T0 = T4 ? T3 : T1;
  assign T1 = T2 ? 5'h0 : v;
  assign T2 = io_enable & io_rst;
  assign T3 = v + 5'h1;
  assign T4 = io_enable & T5;
  assign T5 = io_rst ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      v <= 5'h0;
    end else if(T4) begin
      v <= T3;
    end else if(T2) begin
      v <= 5'h0;
    end
  end
endmodule

module Switch_0(input clk, input reset,
    input  io_signalOn,
    output io_state,
    input  io_rst
);

  wire T0;
  reg  stateReg;
  wire T8;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    stateReg = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_state = T0;
  assign T0 = stateReg | io_signalOn;
  assign T8 = reset ? 1'h0 : T1;
  assign T1 = T6 ? stateReg : T2;
  assign T2 = T4 ? 1'h0 : T3;
  assign T3 = io_signalOn ? 1'h1 : stateReg;
  assign T4 = T5 & io_rst;
  assign T5 = io_signalOn ^ 1'h1;
  assign T6 = T7 ^ 1'h1;
  assign T7 = io_signalOn | io_rst;

  always @(posedge clk) begin
    if(reset) begin
      stateReg <= 1'h0;
    end else if(T6) begin
      stateReg <= stateReg;
    end else if(T4) begin
      stateReg <= 1'h0;
    end else if(io_signalOn) begin
      stateReg <= 1'h1;
    end
  end
endmodule

module Switch_1(input clk, input reset,
    input  io_signalOn,
    output io_state,
    input  io_rst
);

  wire T0;
  reg  stateReg;
  wire T8;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    stateReg = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_state = T0;
  assign T0 = stateReg | io_signalOn;
  assign T8 = reset ? 1'h1 : T1;
  assign T1 = T6 ? stateReg : T2;
  assign T2 = T4 ? 1'h0 : T3;
  assign T3 = io_signalOn ? 1'h1 : stateReg;
  assign T4 = T5 & io_rst;
  assign T5 = io_signalOn ^ 1'h1;
  assign T6 = T7 ^ 1'h1;
  assign T7 = io_signalOn | io_rst;

  always @(posedge clk) begin
    if(reset) begin
      stateReg <= 1'h1;
    end else if(T6) begin
      stateReg <= stateReg;
    end else if(T4) begin
      stateReg <= 1'h0;
    end else if(io_signalOn) begin
      stateReg <= 1'h1;
    end
  end
endmodule

module WarpControl_0(input clk, input reset,
    output io_ready,
    input  io_start,
    input  io_nextReady,
    output io_valid,
    output io_done,
    output[4:0] io_selectX,
    output io_memoryRestart,
    output io_chainRestart
);

  wire signalDone;
  reg  signalTailing;
  wire T8;
  wire signalLastActiveCycle;
  wire signalResetSelectX;
  reg  signalFirstOutputCycle;
  wire T9;
  wire signalOutputtingNext;
  wire T0;
  wire signalFirstReadyCycle;
  wire T1;
  wire signalLastCycleInPass;
  wire signalStartNewPass;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire[5:0] cycleInPass_io_value;
  wire[8:0] cycle_io_value;
  wire[4:0] tailCycle_io_value;
  wire[4:0] selectX_io_value;
  wire isActive_io_state;
  wire isReady_io_state;
  wire isOutputting_io_state;
  wire isTailing_io_state;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    signalTailing = {1{$random}};
    signalFirstOutputCycle = {1{$random}};
  end
// synthesis translate_on
`endif

  assign signalDone = tailCycle_io_value == 5'h1f;
  assign T8 = reset ? 1'h0 : signalLastActiveCycle;
  assign signalLastActiveCycle = cycle_io_value == 9'h187;
  assign signalResetSelectX = selectX_io_value == 5'h1f;
  assign T9 = reset ? 1'h0 : signalOutputtingNext;
  assign signalOutputtingNext = T0 & isActive_io_state;
  assign T0 = cycleInPass_io_value == 6'h30;
  assign signalFirstReadyCycle = T1 & isTailing_io_state;
  assign T1 = tailCycle_io_value == 5'h0;
  assign signalLastCycleInPass = cycleInPass_io_value == 6'h30;
  assign io_chainRestart = signalStartNewPass;
  assign signalStartNewPass = cycleInPass_io_value == 6'h0;
  assign io_memoryRestart = T2;
  assign T2 = T4 & T3;
  assign T3 = io_start ^ 1'h1;
  assign T4 = isReady_io_state | signalLastActiveCycle;
  assign io_selectX = selectX_io_value;
  assign io_done = signalDone;
  assign io_valid = isOutputting_io_state;
  assign io_ready = T5;
  assign T5 = T7 & T6;
  assign T6 = io_start ^ 1'h1;
  assign T7 = isReady_io_state & io_nextReady;
  Counter_0 cycleInPass(.clk(clk), .reset(reset),
       .io_enable( isActive_io_state ),
       .io_rst( signalLastCycleInPass ),
       .io_value( cycleInPass_io_value )
  );
  Counter_3 cycle(.clk(clk), .reset(reset),
       .io_enable( isActive_io_state ),
       .io_rst( signalLastActiveCycle ),
       .io_value( cycle_io_value )
  );
  Counter_4 tailCycle(.clk(clk), .reset(reset),
       .io_enable( isTailing_io_state ),
       .io_rst( signalDone ),
       .io_value( tailCycle_io_value )
  );
  Counter_4 selectX(.clk(clk), .reset(reset),
       .io_enable( isOutputting_io_state ),
       .io_rst( signalResetSelectX ),
       .io_value( selectX_io_value )
  );
  Switch_0 isActive(.clk(clk), .reset(reset),
       .io_signalOn( io_start ),
       .io_state( isActive_io_state ),
       .io_rst( signalLastActiveCycle )
  );
  Switch_1 isReady(.clk(clk), .reset(reset),
       .io_signalOn( signalFirstReadyCycle ),
       .io_state( isReady_io_state ),
       .io_rst( io_start )
  );
  Switch_0 isOutputting(.clk(clk), .reset(reset),
       .io_signalOn( signalFirstOutputCycle ),
       .io_state( isOutputting_io_state ),
       .io_rst( signalResetSelectX )
  );
  Switch_0 isTailing(.clk(clk), .reset(reset),
       .io_signalOn( signalTailing ),
       .io_state( isTailing_io_state ),
       .io_rst( signalDone )
  );

  always @(posedge clk) begin
    if(reset) begin
      signalTailing <= 1'h0;
    end else begin
      signalTailing <= signalLastActiveCycle;
    end
    if(reset) begin
      signalFirstOutputCycle <= 1'h0;
    end else begin
      signalFirstOutputCycle <= signalOutputtingNext;
    end
  end
endmodule

module ProcessingUnit(input clk, input reset,
    input [15:0] io_xs,
    input [15:0] io_ws,
    output[15:0] io_xOut,
    output[9:0] io_yOut,
    input [7:0] io_bias,
    input  io_restartIn,
    output io_restartOut
);

  reg  restartReg;
  wire T54;
  reg [9:0] yReg;
  wire[9:0] T55;
  wire[9:0] T0;
  wire[9:0] T1;
  wire[9:0] T56;
  wire[5:0] T2;
  wire[5:0] T3;
  wire[4:0] innerProd;
  wire[4:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[1:0] T9;
  wire[1:0] T10;
  wire T11;
  wire[15:0] T12;
  wire[15:0] T13;
  wire[1:0] T57;
  wire T14;
  wire[2:0] T58;
  wire[1:0] T15;
  wire[1:0] T16;
  wire T17;
  wire[1:0] T59;
  wire T18;
  wire[3:0] T60;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[1:0] T21;
  wire[1:0] T22;
  wire T23;
  wire[1:0] T61;
  wire T24;
  wire[2:0] T62;
  wire[1:0] T25;
  wire[1:0] T26;
  wire T27;
  wire[1:0] T63;
  wire T28;
  wire[4:0] T64;
  wire[3:0] T29;
  wire[3:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire T35;
  wire[1:0] T65;
  wire T36;
  wire[2:0] T66;
  wire[1:0] T37;
  wire[1:0] T38;
  wire T39;
  wire[1:0] T67;
  wire T40;
  wire[3:0] T68;
  wire[2:0] T41;
  wire[2:0] T42;
  wire[1:0] T43;
  wire[1:0] T44;
  wire T45;
  wire[1:0] T69;
  wire T46;
  wire[2:0] T70;
  wire[1:0] T47;
  wire[1:0] T48;
  wire T49;
  wire[1:0] T71;
  wire T50;
  wire[3:0] T72;
  wire T73;
  wire[9:0] T74;
  wire[7:0] T51;
  wire[7:0] T75;
  wire[5:0] T52;
  wire[5:0] T53;
  wire[1:0] T76;
  wire T77;
  wire[1:0] T78;
  wire T79;
  reg [15:0] xReg;
  wire[15:0] T80;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    restartReg = {1{$random}};
    yReg = {1{$random}};
    xReg = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_restartOut = restartReg;
  assign T54 = reset ? 1'h0 : io_restartIn;
  assign io_yOut = yReg;
  assign T55 = reset ? 10'h0 : T0;
  assign T0 = io_restartIn ? T74 : T1;
  assign T1 = yReg + T56;
  assign T56 = {T72, T2};
  assign T2 = T3;
  assign T3 = {1'h0, innerProd};
  assign innerProd = T64 + T4;
  assign T4 = {1'h0, T5};
  assign T5 = T60 + T6;
  assign T6 = {1'h0, T7};
  assign T7 = T58 + T8;
  assign T8 = {1'h0, T9};
  assign T9 = T57 + T10;
  assign T10 = {1'h0, T11};
  assign T11 = T12[15];
  assign T12 = ~ T13;
  assign T13 = io_xs ^ io_ws;
  assign T57 = {1'h0, T14};
  assign T14 = T12[14];
  assign T58 = {1'h0, T15};
  assign T15 = T59 + T16;
  assign T16 = {1'h0, T17};
  assign T17 = T12[13];
  assign T59 = {1'h0, T18};
  assign T18 = T12[12];
  assign T60 = {1'h0, T19};
  assign T19 = T62 + T20;
  assign T20 = {1'h0, T21};
  assign T21 = T61 + T22;
  assign T22 = {1'h0, T23};
  assign T23 = T12[11];
  assign T61 = {1'h0, T24};
  assign T24 = T12[10];
  assign T62 = {1'h0, T25};
  assign T25 = T63 + T26;
  assign T26 = {1'h0, T27};
  assign T27 = T12[9];
  assign T63 = {1'h0, T28};
  assign T28 = T12[8];
  assign T64 = {1'h0, T29};
  assign T29 = T68 + T30;
  assign T30 = {1'h0, T31};
  assign T31 = T66 + T32;
  assign T32 = {1'h0, T33};
  assign T33 = T65 + T34;
  assign T34 = {1'h0, T35};
  assign T35 = T12[7];
  assign T65 = {1'h0, T36};
  assign T36 = T12[6];
  assign T66 = {1'h0, T37};
  assign T37 = T67 + T38;
  assign T38 = {1'h0, T39};
  assign T39 = T12[5];
  assign T67 = {1'h0, T40};
  assign T40 = T12[4];
  assign T68 = {1'h0, T41};
  assign T41 = T70 + T42;
  assign T42 = {1'h0, T43};
  assign T43 = T69 + T44;
  assign T44 = {1'h0, T45};
  assign T45 = T12[3];
  assign T69 = {1'h0, T46};
  assign T46 = T12[2];
  assign T70 = {1'h0, T47};
  assign T47 = T71 + T48;
  assign T48 = {1'h0, T49};
  assign T49 = T12[1];
  assign T71 = {1'h0, T50};
  assign T50 = T12[0];
  assign T72 = T73 ? 4'hf : 4'h0;
  assign T73 = T2[5];
  assign T74 = {T78, T51};
  assign T51 = io_bias + T75;
  assign T75 = {T76, T52};
  assign T52 = T53;
  assign T53 = {1'h0, innerProd};
  assign T76 = T77 ? 2'h3 : 2'h0;
  assign T77 = T52[5];
  assign T78 = T79 ? 2'h3 : 2'h0;
  assign T79 = T51[7];
  assign io_xOut = xReg;
  assign T80 = reset ? 16'h0 : io_xs;

  always @(posedge clk) begin
    if(reset) begin
      restartReg <= 1'h0;
    end else begin
      restartReg <= io_restartIn;
    end
    if(reset) begin
      yReg <= 10'h0;
    end else if(io_restartIn) begin
      yReg <= T74;
    end else begin
      yReg <= T1;
    end
    if(reset) begin
      xReg <= 16'h0;
    end else begin
      xReg <= io_xs;
    end
  end
endmodule

module Chain_0(input clk, input reset,
    input [15:0] io_weights_31,
    input [15:0] io_weights_30,
    input [15:0] io_weights_29,
    input [15:0] io_weights_28,
    input [15:0] io_weights_27,
    input [15:0] io_weights_26,
    input [15:0] io_weights_25,
    input [15:0] io_weights_24,
    input [15:0] io_weights_23,
    input [15:0] io_weights_22,
    input [15:0] io_weights_21,
    input [15:0] io_weights_20,
    input [15:0] io_weights_19,
    input [15:0] io_weights_18,
    input [15:0] io_weights_17,
    input [15:0] io_weights_16,
    input [15:0] io_weights_15,
    input [15:0] io_weights_14,
    input [15:0] io_weights_13,
    input [15:0] io_weights_12,
    input [15:0] io_weights_11,
    input [15:0] io_weights_10,
    input [15:0] io_weights_9,
    input [15:0] io_weights_8,
    input [15:0] io_weights_7,
    input [15:0] io_weights_6,
    input [15:0] io_weights_5,
    input [15:0] io_weights_4,
    input [15:0] io_weights_3,
    input [15:0] io_weights_2,
    input [15:0] io_weights_1,
    input [15:0] io_weights_0,
    input [7:0] io_bias,
    input  io_restartIn,
    input [15:0] io_xs,
    output[9:0] io_ys_31,
    output[9:0] io_ys_30,
    output[9:0] io_ys_29,
    output[9:0] io_ys_28,
    output[9:0] io_ys_27,
    output[9:0] io_ys_26,
    output[9:0] io_ys_25,
    output[9:0] io_ys_24,
    output[9:0] io_ys_23,
    output[9:0] io_ys_22,
    output[9:0] io_ys_21,
    output[9:0] io_ys_20,
    output[9:0] io_ys_19,
    output[9:0] io_ys_18,
    output[9:0] io_ys_17,
    output[9:0] io_ys_16,
    output[9:0] io_ys_15,
    output[9:0] io_ys_14,
    output[9:0] io_ys_13,
    output[9:0] io_ys_12,
    output[9:0] io_ys_11,
    output[9:0] io_ys_10,
    output[9:0] io_ys_9,
    output[9:0] io_ys_8,
    output[9:0] io_ys_7,
    output[9:0] io_ys_6,
    output[9:0] io_ys_5,
    output[9:0] io_ys_4,
    output[9:0] io_ys_3,
    output[9:0] io_ys_2,
    output[9:0] io_ys_1,
    output[9:0] io_ys_0
);

  wire[7:0] T64;
  wire[8:0] T0;
  wire[8:0] T1;
  wire[7:0] T65;
  wire[8:0] T2;
  wire[8:0] T3;
  wire[7:0] T66;
  wire[8:0] T4;
  wire[8:0] T5;
  wire[7:0] T67;
  wire[8:0] T6;
  wire[8:0] T7;
  wire[7:0] T68;
  wire[8:0] T8;
  wire[8:0] T9;
  wire[7:0] T69;
  wire[8:0] T10;
  wire[8:0] T11;
  wire[7:0] T70;
  wire[8:0] T12;
  wire[8:0] T13;
  wire[7:0] T71;
  wire[8:0] T14;
  wire[8:0] T15;
  wire[7:0] T72;
  wire[8:0] T16;
  wire[8:0] T17;
  wire[7:0] T73;
  wire[8:0] T18;
  wire[8:0] T19;
  wire[7:0] T74;
  wire[8:0] T20;
  wire[8:0] T21;
  wire[7:0] T75;
  wire[8:0] T22;
  wire[8:0] T23;
  wire[7:0] T76;
  wire[8:0] T24;
  wire[8:0] T25;
  wire[7:0] T77;
  wire[8:0] T26;
  wire[8:0] T27;
  wire[7:0] T78;
  wire[8:0] T28;
  wire[8:0] T29;
  wire[7:0] T79;
  wire[8:0] T30;
  wire[8:0] T31;
  wire[7:0] T80;
  wire[8:0] T32;
  wire[8:0] T33;
  wire[7:0] T81;
  wire[8:0] T34;
  wire[8:0] T35;
  wire[7:0] T82;
  wire[8:0] T36;
  wire[8:0] T37;
  wire[7:0] T83;
  wire[8:0] T38;
  wire[8:0] T39;
  wire[7:0] T84;
  wire[8:0] T40;
  wire[8:0] T41;
  wire[7:0] T85;
  wire[8:0] T42;
  wire[8:0] T43;
  wire[7:0] T86;
  wire[8:0] T44;
  wire[8:0] T45;
  wire[7:0] T87;
  wire[8:0] T46;
  wire[8:0] T47;
  wire[7:0] T88;
  wire[8:0] T48;
  wire[8:0] T49;
  wire[7:0] T89;
  wire[8:0] T50;
  wire[8:0] T51;
  wire[7:0] T90;
  wire[8:0] T52;
  wire[8:0] T53;
  wire[7:0] T91;
  wire[8:0] T54;
  wire[8:0] T55;
  wire[7:0] T92;
  wire[8:0] T56;
  wire[8:0] T57;
  wire[7:0] T93;
  wire[8:0] T58;
  wire[8:0] T59;
  wire[7:0] T94;
  wire[8:0] T60;
  wire[8:0] T61;
  wire[7:0] T95;
  wire[8:0] T62;
  wire[8:0] T63;
  wire[15:0] ProcessingUnit_io_xOut;
  wire[9:0] ProcessingUnit_io_yOut;
  wire ProcessingUnit_io_restartOut;
  wire[15:0] ProcessingUnit_1_io_xOut;
  wire[9:0] ProcessingUnit_1_io_yOut;
  wire ProcessingUnit_1_io_restartOut;
  wire[15:0] ProcessingUnit_2_io_xOut;
  wire[9:0] ProcessingUnit_2_io_yOut;
  wire ProcessingUnit_2_io_restartOut;
  wire[15:0] ProcessingUnit_3_io_xOut;
  wire[9:0] ProcessingUnit_3_io_yOut;
  wire ProcessingUnit_3_io_restartOut;
  wire[15:0] ProcessingUnit_4_io_xOut;
  wire[9:0] ProcessingUnit_4_io_yOut;
  wire ProcessingUnit_4_io_restartOut;
  wire[15:0] ProcessingUnit_5_io_xOut;
  wire[9:0] ProcessingUnit_5_io_yOut;
  wire ProcessingUnit_5_io_restartOut;
  wire[15:0] ProcessingUnit_6_io_xOut;
  wire[9:0] ProcessingUnit_6_io_yOut;
  wire ProcessingUnit_6_io_restartOut;
  wire[15:0] ProcessingUnit_7_io_xOut;
  wire[9:0] ProcessingUnit_7_io_yOut;
  wire ProcessingUnit_7_io_restartOut;
  wire[15:0] ProcessingUnit_8_io_xOut;
  wire[9:0] ProcessingUnit_8_io_yOut;
  wire ProcessingUnit_8_io_restartOut;
  wire[15:0] ProcessingUnit_9_io_xOut;
  wire[9:0] ProcessingUnit_9_io_yOut;
  wire ProcessingUnit_9_io_restartOut;
  wire[15:0] ProcessingUnit_10_io_xOut;
  wire[9:0] ProcessingUnit_10_io_yOut;
  wire ProcessingUnit_10_io_restartOut;
  wire[15:0] ProcessingUnit_11_io_xOut;
  wire[9:0] ProcessingUnit_11_io_yOut;
  wire ProcessingUnit_11_io_restartOut;
  wire[15:0] ProcessingUnit_12_io_xOut;
  wire[9:0] ProcessingUnit_12_io_yOut;
  wire ProcessingUnit_12_io_restartOut;
  wire[15:0] ProcessingUnit_13_io_xOut;
  wire[9:0] ProcessingUnit_13_io_yOut;
  wire ProcessingUnit_13_io_restartOut;
  wire[15:0] ProcessingUnit_14_io_xOut;
  wire[9:0] ProcessingUnit_14_io_yOut;
  wire ProcessingUnit_14_io_restartOut;
  wire[15:0] ProcessingUnit_15_io_xOut;
  wire[9:0] ProcessingUnit_15_io_yOut;
  wire ProcessingUnit_15_io_restartOut;
  wire[15:0] ProcessingUnit_16_io_xOut;
  wire[9:0] ProcessingUnit_16_io_yOut;
  wire ProcessingUnit_16_io_restartOut;
  wire[15:0] ProcessingUnit_17_io_xOut;
  wire[9:0] ProcessingUnit_17_io_yOut;
  wire ProcessingUnit_17_io_restartOut;
  wire[15:0] ProcessingUnit_18_io_xOut;
  wire[9:0] ProcessingUnit_18_io_yOut;
  wire ProcessingUnit_18_io_restartOut;
  wire[15:0] ProcessingUnit_19_io_xOut;
  wire[9:0] ProcessingUnit_19_io_yOut;
  wire ProcessingUnit_19_io_restartOut;
  wire[15:0] ProcessingUnit_20_io_xOut;
  wire[9:0] ProcessingUnit_20_io_yOut;
  wire ProcessingUnit_20_io_restartOut;
  wire[15:0] ProcessingUnit_21_io_xOut;
  wire[9:0] ProcessingUnit_21_io_yOut;
  wire ProcessingUnit_21_io_restartOut;
  wire[15:0] ProcessingUnit_22_io_xOut;
  wire[9:0] ProcessingUnit_22_io_yOut;
  wire ProcessingUnit_22_io_restartOut;
  wire[15:0] ProcessingUnit_23_io_xOut;
  wire[9:0] ProcessingUnit_23_io_yOut;
  wire ProcessingUnit_23_io_restartOut;
  wire[15:0] ProcessingUnit_24_io_xOut;
  wire[9:0] ProcessingUnit_24_io_yOut;
  wire ProcessingUnit_24_io_restartOut;
  wire[15:0] ProcessingUnit_25_io_xOut;
  wire[9:0] ProcessingUnit_25_io_yOut;
  wire ProcessingUnit_25_io_restartOut;
  wire[15:0] ProcessingUnit_26_io_xOut;
  wire[9:0] ProcessingUnit_26_io_yOut;
  wire ProcessingUnit_26_io_restartOut;
  wire[15:0] ProcessingUnit_27_io_xOut;
  wire[9:0] ProcessingUnit_27_io_yOut;
  wire ProcessingUnit_27_io_restartOut;
  wire[15:0] ProcessingUnit_28_io_xOut;
  wire[9:0] ProcessingUnit_28_io_yOut;
  wire ProcessingUnit_28_io_restartOut;
  wire[15:0] ProcessingUnit_29_io_xOut;
  wire[9:0] ProcessingUnit_29_io_yOut;
  wire ProcessingUnit_29_io_restartOut;
  wire[15:0] ProcessingUnit_30_io_xOut;
  wire[9:0] ProcessingUnit_30_io_yOut;
  wire ProcessingUnit_30_io_restartOut;
  wire[9:0] ProcessingUnit_31_io_yOut;


  assign T64 = T0[7:0];
  assign T0 = T1;
  assign T1 = {1'h0, io_bias};
  assign T65 = T2[7:0];
  assign T2 = T3;
  assign T3 = {1'h0, io_bias};
  assign T66 = T4[7:0];
  assign T4 = T5;
  assign T5 = {1'h0, io_bias};
  assign T67 = T6[7:0];
  assign T6 = T7;
  assign T7 = {1'h0, io_bias};
  assign T68 = T8[7:0];
  assign T8 = T9;
  assign T9 = {1'h0, io_bias};
  assign T69 = T10[7:0];
  assign T10 = T11;
  assign T11 = {1'h0, io_bias};
  assign T70 = T12[7:0];
  assign T12 = T13;
  assign T13 = {1'h0, io_bias};
  assign T71 = T14[7:0];
  assign T14 = T15;
  assign T15 = {1'h0, io_bias};
  assign T72 = T16[7:0];
  assign T16 = T17;
  assign T17 = {1'h0, io_bias};
  assign T73 = T18[7:0];
  assign T18 = T19;
  assign T19 = {1'h0, io_bias};
  assign T74 = T20[7:0];
  assign T20 = T21;
  assign T21 = {1'h0, io_bias};
  assign T75 = T22[7:0];
  assign T22 = T23;
  assign T23 = {1'h0, io_bias};
  assign T76 = T24[7:0];
  assign T24 = T25;
  assign T25 = {1'h0, io_bias};
  assign T77 = T26[7:0];
  assign T26 = T27;
  assign T27 = {1'h0, io_bias};
  assign T78 = T28[7:0];
  assign T28 = T29;
  assign T29 = {1'h0, io_bias};
  assign T79 = T30[7:0];
  assign T30 = T31;
  assign T31 = {1'h0, io_bias};
  assign T80 = T32[7:0];
  assign T32 = T33;
  assign T33 = {1'h0, io_bias};
  assign T81 = T34[7:0];
  assign T34 = T35;
  assign T35 = {1'h0, io_bias};
  assign T82 = T36[7:0];
  assign T36 = T37;
  assign T37 = {1'h0, io_bias};
  assign T83 = T38[7:0];
  assign T38 = T39;
  assign T39 = {1'h0, io_bias};
  assign T84 = T40[7:0];
  assign T40 = T41;
  assign T41 = {1'h0, io_bias};
  assign T85 = T42[7:0];
  assign T42 = T43;
  assign T43 = {1'h0, io_bias};
  assign T86 = T44[7:0];
  assign T44 = T45;
  assign T45 = {1'h0, io_bias};
  assign T87 = T46[7:0];
  assign T46 = T47;
  assign T47 = {1'h0, io_bias};
  assign T88 = T48[7:0];
  assign T48 = T49;
  assign T49 = {1'h0, io_bias};
  assign T89 = T50[7:0];
  assign T50 = T51;
  assign T51 = {1'h0, io_bias};
  assign T90 = T52[7:0];
  assign T52 = T53;
  assign T53 = {1'h0, io_bias};
  assign T91 = T54[7:0];
  assign T54 = T55;
  assign T55 = {1'h0, io_bias};
  assign T92 = T56[7:0];
  assign T56 = T57;
  assign T57 = {1'h0, io_bias};
  assign T93 = T58[7:0];
  assign T58 = T59;
  assign T59 = {1'h0, io_bias};
  assign T94 = T60[7:0];
  assign T60 = T61;
  assign T61 = {1'h0, io_bias};
  assign T95 = T62[7:0];
  assign T62 = T63;
  assign T63 = {1'h0, io_bias};
  assign io_ys_0 = ProcessingUnit_io_yOut;
  assign io_ys_1 = ProcessingUnit_1_io_yOut;
  assign io_ys_2 = ProcessingUnit_2_io_yOut;
  assign io_ys_3 = ProcessingUnit_3_io_yOut;
  assign io_ys_4 = ProcessingUnit_4_io_yOut;
  assign io_ys_5 = ProcessingUnit_5_io_yOut;
  assign io_ys_6 = ProcessingUnit_6_io_yOut;
  assign io_ys_7 = ProcessingUnit_7_io_yOut;
  assign io_ys_8 = ProcessingUnit_8_io_yOut;
  assign io_ys_9 = ProcessingUnit_9_io_yOut;
  assign io_ys_10 = ProcessingUnit_10_io_yOut;
  assign io_ys_11 = ProcessingUnit_11_io_yOut;
  assign io_ys_12 = ProcessingUnit_12_io_yOut;
  assign io_ys_13 = ProcessingUnit_13_io_yOut;
  assign io_ys_14 = ProcessingUnit_14_io_yOut;
  assign io_ys_15 = ProcessingUnit_15_io_yOut;
  assign io_ys_16 = ProcessingUnit_16_io_yOut;
  assign io_ys_17 = ProcessingUnit_17_io_yOut;
  assign io_ys_18 = ProcessingUnit_18_io_yOut;
  assign io_ys_19 = ProcessingUnit_19_io_yOut;
  assign io_ys_20 = ProcessingUnit_20_io_yOut;
  assign io_ys_21 = ProcessingUnit_21_io_yOut;
  assign io_ys_22 = ProcessingUnit_22_io_yOut;
  assign io_ys_23 = ProcessingUnit_23_io_yOut;
  assign io_ys_24 = ProcessingUnit_24_io_yOut;
  assign io_ys_25 = ProcessingUnit_25_io_yOut;
  assign io_ys_26 = ProcessingUnit_26_io_yOut;
  assign io_ys_27 = ProcessingUnit_27_io_yOut;
  assign io_ys_28 = ProcessingUnit_28_io_yOut;
  assign io_ys_29 = ProcessingUnit_29_io_yOut;
  assign io_ys_30 = ProcessingUnit_30_io_yOut;
  assign io_ys_31 = ProcessingUnit_31_io_yOut;
  ProcessingUnit ProcessingUnit(.clk(clk), .reset(reset),
       .io_xs( io_xs ),
       .io_ws( io_weights_0 ),
       .io_xOut( ProcessingUnit_io_xOut ),
       .io_yOut( ProcessingUnit_io_yOut ),
       .io_bias( T95 ),
       .io_restartIn( io_restartIn ),
       .io_restartOut( ProcessingUnit_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_1(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_io_xOut ),
       .io_ws( io_weights_1 ),
       .io_xOut( ProcessingUnit_1_io_xOut ),
       .io_yOut( ProcessingUnit_1_io_yOut ),
       .io_bias( T94 ),
       .io_restartIn( ProcessingUnit_io_restartOut ),
       .io_restartOut( ProcessingUnit_1_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_2(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_1_io_xOut ),
       .io_ws( io_weights_2 ),
       .io_xOut( ProcessingUnit_2_io_xOut ),
       .io_yOut( ProcessingUnit_2_io_yOut ),
       .io_bias( T93 ),
       .io_restartIn( ProcessingUnit_1_io_restartOut ),
       .io_restartOut( ProcessingUnit_2_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_3(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_2_io_xOut ),
       .io_ws( io_weights_3 ),
       .io_xOut( ProcessingUnit_3_io_xOut ),
       .io_yOut( ProcessingUnit_3_io_yOut ),
       .io_bias( T92 ),
       .io_restartIn( ProcessingUnit_2_io_restartOut ),
       .io_restartOut( ProcessingUnit_3_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_4(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_3_io_xOut ),
       .io_ws( io_weights_4 ),
       .io_xOut( ProcessingUnit_4_io_xOut ),
       .io_yOut( ProcessingUnit_4_io_yOut ),
       .io_bias( T91 ),
       .io_restartIn( ProcessingUnit_3_io_restartOut ),
       .io_restartOut( ProcessingUnit_4_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_5(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_4_io_xOut ),
       .io_ws( io_weights_5 ),
       .io_xOut( ProcessingUnit_5_io_xOut ),
       .io_yOut( ProcessingUnit_5_io_yOut ),
       .io_bias( T90 ),
       .io_restartIn( ProcessingUnit_4_io_restartOut ),
       .io_restartOut( ProcessingUnit_5_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_6(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_5_io_xOut ),
       .io_ws( io_weights_6 ),
       .io_xOut( ProcessingUnit_6_io_xOut ),
       .io_yOut( ProcessingUnit_6_io_yOut ),
       .io_bias( T89 ),
       .io_restartIn( ProcessingUnit_5_io_restartOut ),
       .io_restartOut( ProcessingUnit_6_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_7(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_6_io_xOut ),
       .io_ws( io_weights_7 ),
       .io_xOut( ProcessingUnit_7_io_xOut ),
       .io_yOut( ProcessingUnit_7_io_yOut ),
       .io_bias( T88 ),
       .io_restartIn( ProcessingUnit_6_io_restartOut ),
       .io_restartOut( ProcessingUnit_7_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_8(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_7_io_xOut ),
       .io_ws( io_weights_8 ),
       .io_xOut( ProcessingUnit_8_io_xOut ),
       .io_yOut( ProcessingUnit_8_io_yOut ),
       .io_bias( T87 ),
       .io_restartIn( ProcessingUnit_7_io_restartOut ),
       .io_restartOut( ProcessingUnit_8_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_9(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_8_io_xOut ),
       .io_ws( io_weights_9 ),
       .io_xOut( ProcessingUnit_9_io_xOut ),
       .io_yOut( ProcessingUnit_9_io_yOut ),
       .io_bias( T86 ),
       .io_restartIn( ProcessingUnit_8_io_restartOut ),
       .io_restartOut( ProcessingUnit_9_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_10(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_9_io_xOut ),
       .io_ws( io_weights_10 ),
       .io_xOut( ProcessingUnit_10_io_xOut ),
       .io_yOut( ProcessingUnit_10_io_yOut ),
       .io_bias( T85 ),
       .io_restartIn( ProcessingUnit_9_io_restartOut ),
       .io_restartOut( ProcessingUnit_10_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_11(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_10_io_xOut ),
       .io_ws( io_weights_11 ),
       .io_xOut( ProcessingUnit_11_io_xOut ),
       .io_yOut( ProcessingUnit_11_io_yOut ),
       .io_bias( T84 ),
       .io_restartIn( ProcessingUnit_10_io_restartOut ),
       .io_restartOut( ProcessingUnit_11_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_12(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_11_io_xOut ),
       .io_ws( io_weights_12 ),
       .io_xOut( ProcessingUnit_12_io_xOut ),
       .io_yOut( ProcessingUnit_12_io_yOut ),
       .io_bias( T83 ),
       .io_restartIn( ProcessingUnit_11_io_restartOut ),
       .io_restartOut( ProcessingUnit_12_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_13(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_12_io_xOut ),
       .io_ws( io_weights_13 ),
       .io_xOut( ProcessingUnit_13_io_xOut ),
       .io_yOut( ProcessingUnit_13_io_yOut ),
       .io_bias( T82 ),
       .io_restartIn( ProcessingUnit_12_io_restartOut ),
       .io_restartOut( ProcessingUnit_13_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_14(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_13_io_xOut ),
       .io_ws( io_weights_14 ),
       .io_xOut( ProcessingUnit_14_io_xOut ),
       .io_yOut( ProcessingUnit_14_io_yOut ),
       .io_bias( T81 ),
       .io_restartIn( ProcessingUnit_13_io_restartOut ),
       .io_restartOut( ProcessingUnit_14_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_15(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_14_io_xOut ),
       .io_ws( io_weights_15 ),
       .io_xOut( ProcessingUnit_15_io_xOut ),
       .io_yOut( ProcessingUnit_15_io_yOut ),
       .io_bias( T80 ),
       .io_restartIn( ProcessingUnit_14_io_restartOut ),
       .io_restartOut( ProcessingUnit_15_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_16(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_15_io_xOut ),
       .io_ws( io_weights_16 ),
       .io_xOut( ProcessingUnit_16_io_xOut ),
       .io_yOut( ProcessingUnit_16_io_yOut ),
       .io_bias( T79 ),
       .io_restartIn( ProcessingUnit_15_io_restartOut ),
       .io_restartOut( ProcessingUnit_16_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_17(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_16_io_xOut ),
       .io_ws( io_weights_17 ),
       .io_xOut( ProcessingUnit_17_io_xOut ),
       .io_yOut( ProcessingUnit_17_io_yOut ),
       .io_bias( T78 ),
       .io_restartIn( ProcessingUnit_16_io_restartOut ),
       .io_restartOut( ProcessingUnit_17_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_18(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_17_io_xOut ),
       .io_ws( io_weights_18 ),
       .io_xOut( ProcessingUnit_18_io_xOut ),
       .io_yOut( ProcessingUnit_18_io_yOut ),
       .io_bias( T77 ),
       .io_restartIn( ProcessingUnit_17_io_restartOut ),
       .io_restartOut( ProcessingUnit_18_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_19(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_18_io_xOut ),
       .io_ws( io_weights_19 ),
       .io_xOut( ProcessingUnit_19_io_xOut ),
       .io_yOut( ProcessingUnit_19_io_yOut ),
       .io_bias( T76 ),
       .io_restartIn( ProcessingUnit_18_io_restartOut ),
       .io_restartOut( ProcessingUnit_19_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_20(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_19_io_xOut ),
       .io_ws( io_weights_20 ),
       .io_xOut( ProcessingUnit_20_io_xOut ),
       .io_yOut( ProcessingUnit_20_io_yOut ),
       .io_bias( T75 ),
       .io_restartIn( ProcessingUnit_19_io_restartOut ),
       .io_restartOut( ProcessingUnit_20_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_21(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_20_io_xOut ),
       .io_ws( io_weights_21 ),
       .io_xOut( ProcessingUnit_21_io_xOut ),
       .io_yOut( ProcessingUnit_21_io_yOut ),
       .io_bias( T74 ),
       .io_restartIn( ProcessingUnit_20_io_restartOut ),
       .io_restartOut( ProcessingUnit_21_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_22(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_21_io_xOut ),
       .io_ws( io_weights_22 ),
       .io_xOut( ProcessingUnit_22_io_xOut ),
       .io_yOut( ProcessingUnit_22_io_yOut ),
       .io_bias( T73 ),
       .io_restartIn( ProcessingUnit_21_io_restartOut ),
       .io_restartOut( ProcessingUnit_22_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_23(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_22_io_xOut ),
       .io_ws( io_weights_23 ),
       .io_xOut( ProcessingUnit_23_io_xOut ),
       .io_yOut( ProcessingUnit_23_io_yOut ),
       .io_bias( T72 ),
       .io_restartIn( ProcessingUnit_22_io_restartOut ),
       .io_restartOut( ProcessingUnit_23_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_24(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_23_io_xOut ),
       .io_ws( io_weights_24 ),
       .io_xOut( ProcessingUnit_24_io_xOut ),
       .io_yOut( ProcessingUnit_24_io_yOut ),
       .io_bias( T71 ),
       .io_restartIn( ProcessingUnit_23_io_restartOut ),
       .io_restartOut( ProcessingUnit_24_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_25(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_24_io_xOut ),
       .io_ws( io_weights_25 ),
       .io_xOut( ProcessingUnit_25_io_xOut ),
       .io_yOut( ProcessingUnit_25_io_yOut ),
       .io_bias( T70 ),
       .io_restartIn( ProcessingUnit_24_io_restartOut ),
       .io_restartOut( ProcessingUnit_25_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_26(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_25_io_xOut ),
       .io_ws( io_weights_26 ),
       .io_xOut( ProcessingUnit_26_io_xOut ),
       .io_yOut( ProcessingUnit_26_io_yOut ),
       .io_bias( T69 ),
       .io_restartIn( ProcessingUnit_25_io_restartOut ),
       .io_restartOut( ProcessingUnit_26_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_27(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_26_io_xOut ),
       .io_ws( io_weights_27 ),
       .io_xOut( ProcessingUnit_27_io_xOut ),
       .io_yOut( ProcessingUnit_27_io_yOut ),
       .io_bias( T68 ),
       .io_restartIn( ProcessingUnit_26_io_restartOut ),
       .io_restartOut( ProcessingUnit_27_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_28(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_27_io_xOut ),
       .io_ws( io_weights_28 ),
       .io_xOut( ProcessingUnit_28_io_xOut ),
       .io_yOut( ProcessingUnit_28_io_yOut ),
       .io_bias( T67 ),
       .io_restartIn( ProcessingUnit_27_io_restartOut ),
       .io_restartOut( ProcessingUnit_28_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_29(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_28_io_xOut ),
       .io_ws( io_weights_29 ),
       .io_xOut( ProcessingUnit_29_io_xOut ),
       .io_yOut( ProcessingUnit_29_io_yOut ),
       .io_bias( T66 ),
       .io_restartIn( ProcessingUnit_28_io_restartOut ),
       .io_restartOut( ProcessingUnit_29_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_30(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_29_io_xOut ),
       .io_ws( io_weights_30 ),
       .io_xOut( ProcessingUnit_30_io_xOut ),
       .io_yOut( ProcessingUnit_30_io_yOut ),
       .io_bias( T65 ),
       .io_restartIn( ProcessingUnit_29_io_restartOut ),
       .io_restartOut( ProcessingUnit_30_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_31(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_30_io_xOut ),
       .io_ws( io_weights_31 ),
       //.io_xOut(  )
       .io_yOut( ProcessingUnit_31_io_yOut ),
       .io_bias( T64 ),
       .io_restartIn( ProcessingUnit_30_io_restartOut )
       //.io_restartOut(  )
  );
endmodule

module Activation_0(
    input [9:0] io_in_31,
    input [9:0] io_in_30,
    input [9:0] io_in_29,
    input [9:0] io_in_28,
    input [9:0] io_in_27,
    input [9:0] io_in_26,
    input [9:0] io_in_25,
    input [9:0] io_in_24,
    input [9:0] io_in_23,
    input [9:0] io_in_22,
    input [9:0] io_in_21,
    input [9:0] io_in_20,
    input [9:0] io_in_19,
    input [9:0] io_in_18,
    input [9:0] io_in_17,
    input [9:0] io_in_16,
    input [9:0] io_in_15,
    input [9:0] io_in_14,
    input [9:0] io_in_13,
    input [9:0] io_in_12,
    input [9:0] io_in_11,
    input [9:0] io_in_10,
    input [9:0] io_in_9,
    input [9:0] io_in_8,
    input [9:0] io_in_7,
    input [9:0] io_in_6,
    input [9:0] io_in_5,
    input [9:0] io_in_4,
    input [9:0] io_in_3,
    input [9:0] io_in_2,
    input [9:0] io_in_1,
    input [9:0] io_in_0,
    output io_out_31,
    output io_out_30,
    output io_out_29,
    output io_out_28,
    output io_out_27,
    output io_out_26,
    output io_out_25,
    output io_out_24,
    output io_out_23,
    output io_out_22,
    output io_out_21,
    output io_out_20,
    output io_out_19,
    output io_out_18,
    output io_out_17,
    output io_out_16,
    output io_out_15,
    output io_out_14,
    output io_out_13,
    output io_out_12,
    output io_out_11,
    output io_out_10,
    output io_out_9,
    output io_out_8,
    output io_out_7,
    output io_out_6,
    output io_out_5,
    output io_out_4,
    output io_out_3,
    output io_out_2,
    output io_out_1,
    output io_out_0
);

  wire T0;
  wire T1;
  wire[12:0] T2;
  wire[12:0] T3;
  wire T4;
  wire T5;
  wire[12:0] T6;
  wire[12:0] T7;
  wire T8;
  wire T9;
  wire[12:0] T10;
  wire[12:0] T11;
  wire T12;
  wire T13;
  wire[12:0] T14;
  wire[12:0] T15;
  wire T16;
  wire T17;
  wire[12:0] T18;
  wire[12:0] T19;
  wire T20;
  wire T21;
  wire[12:0] T22;
  wire[12:0] T23;
  wire T24;
  wire T25;
  wire[12:0] T26;
  wire[12:0] T27;
  wire T28;
  wire T29;
  wire[12:0] T30;
  wire[12:0] T31;
  wire T32;
  wire T33;
  wire[12:0] T34;
  wire[12:0] T35;
  wire T36;
  wire T37;
  wire[12:0] T38;
  wire[12:0] T39;
  wire T40;
  wire T41;
  wire[12:0] T42;
  wire[12:0] T43;
  wire T44;
  wire T45;
  wire[12:0] T46;
  wire[12:0] T47;
  wire T48;
  wire T49;
  wire[12:0] T50;
  wire[12:0] T51;
  wire T52;
  wire T53;
  wire[12:0] T54;
  wire[12:0] T55;
  wire T56;
  wire T57;
  wire[12:0] T58;
  wire[12:0] T59;
  wire T60;
  wire T61;
  wire[12:0] T62;
  wire[12:0] T63;
  wire T64;
  wire T65;
  wire[12:0] T66;
  wire[12:0] T67;
  wire T68;
  wire T69;
  wire[12:0] T70;
  wire[12:0] T71;
  wire T72;
  wire T73;
  wire[12:0] T74;
  wire[12:0] T75;
  wire T76;
  wire T77;
  wire[12:0] T78;
  wire[12:0] T79;
  wire T80;
  wire T81;
  wire[12:0] T82;
  wire[12:0] T83;
  wire T84;
  wire T85;
  wire[12:0] T86;
  wire[12:0] T87;
  wire T88;
  wire T89;
  wire[12:0] T90;
  wire[12:0] T91;
  wire T92;
  wire T93;
  wire[12:0] T94;
  wire[12:0] T95;
  wire T96;
  wire T97;
  wire[12:0] T98;
  wire[12:0] T99;
  wire T100;
  wire T101;
  wire[12:0] T102;
  wire[12:0] T103;
  wire T104;
  wire T105;
  wire[12:0] T106;
  wire[12:0] T107;
  wire T108;
  wire T109;
  wire[12:0] T110;
  wire[12:0] T111;
  wire T112;
  wire T113;
  wire[12:0] T114;
  wire[12:0] T115;
  wire T116;
  wire T117;
  wire[12:0] T118;
  wire[12:0] T119;
  wire T120;
  wire T121;
  wire[12:0] T122;
  wire[12:0] T123;
  wire T124;
  wire T125;
  wire[12:0] T126;
  wire[12:0] T127;


  assign io_out_0 = T0;
  assign T0 = ~ T1;
  assign T1 = T2[9];
  assign T2 = T3 - 13'h310;
  assign T3 = $signed(io_in_0) * $signed(3'h2);
  assign io_out_1 = T4;
  assign T4 = ~ T5;
  assign T5 = T6[9];
  assign T6 = T7 - 13'h310;
  assign T7 = $signed(io_in_1) * $signed(3'h2);
  assign io_out_2 = T8;
  assign T8 = ~ T9;
  assign T9 = T10[9];
  assign T10 = T11 - 13'h310;
  assign T11 = $signed(io_in_2) * $signed(3'h2);
  assign io_out_3 = T12;
  assign T12 = ~ T13;
  assign T13 = T14[9];
  assign T14 = T15 - 13'h310;
  assign T15 = $signed(io_in_3) * $signed(3'h2);
  assign io_out_4 = T16;
  assign T16 = ~ T17;
  assign T17 = T18[9];
  assign T18 = T19 - 13'h310;
  assign T19 = $signed(io_in_4) * $signed(3'h2);
  assign io_out_5 = T20;
  assign T20 = ~ T21;
  assign T21 = T22[9];
  assign T22 = T23 - 13'h310;
  assign T23 = $signed(io_in_5) * $signed(3'h2);
  assign io_out_6 = T24;
  assign T24 = ~ T25;
  assign T25 = T26[9];
  assign T26 = T27 - 13'h310;
  assign T27 = $signed(io_in_6) * $signed(3'h2);
  assign io_out_7 = T28;
  assign T28 = ~ T29;
  assign T29 = T30[9];
  assign T30 = T31 - 13'h310;
  assign T31 = $signed(io_in_7) * $signed(3'h2);
  assign io_out_8 = T32;
  assign T32 = ~ T33;
  assign T33 = T34[9];
  assign T34 = T35 - 13'h310;
  assign T35 = $signed(io_in_8) * $signed(3'h2);
  assign io_out_9 = T36;
  assign T36 = ~ T37;
  assign T37 = T38[9];
  assign T38 = T39 - 13'h310;
  assign T39 = $signed(io_in_9) * $signed(3'h2);
  assign io_out_10 = T40;
  assign T40 = ~ T41;
  assign T41 = T42[9];
  assign T42 = T43 - 13'h310;
  assign T43 = $signed(io_in_10) * $signed(3'h2);
  assign io_out_11 = T44;
  assign T44 = ~ T45;
  assign T45 = T46[9];
  assign T46 = T47 - 13'h310;
  assign T47 = $signed(io_in_11) * $signed(3'h2);
  assign io_out_12 = T48;
  assign T48 = ~ T49;
  assign T49 = T50[9];
  assign T50 = T51 - 13'h310;
  assign T51 = $signed(io_in_12) * $signed(3'h2);
  assign io_out_13 = T52;
  assign T52 = ~ T53;
  assign T53 = T54[9];
  assign T54 = T55 - 13'h310;
  assign T55 = $signed(io_in_13) * $signed(3'h2);
  assign io_out_14 = T56;
  assign T56 = ~ T57;
  assign T57 = T58[9];
  assign T58 = T59 - 13'h310;
  assign T59 = $signed(io_in_14) * $signed(3'h2);
  assign io_out_15 = T60;
  assign T60 = ~ T61;
  assign T61 = T62[9];
  assign T62 = T63 - 13'h310;
  assign T63 = $signed(io_in_15) * $signed(3'h2);
  assign io_out_16 = T64;
  assign T64 = ~ T65;
  assign T65 = T66[9];
  assign T66 = T67 - 13'h310;
  assign T67 = $signed(io_in_16) * $signed(3'h2);
  assign io_out_17 = T68;
  assign T68 = ~ T69;
  assign T69 = T70[9];
  assign T70 = T71 - 13'h310;
  assign T71 = $signed(io_in_17) * $signed(3'h2);
  assign io_out_18 = T72;
  assign T72 = ~ T73;
  assign T73 = T74[9];
  assign T74 = T75 - 13'h310;
  assign T75 = $signed(io_in_18) * $signed(3'h2);
  assign io_out_19 = T76;
  assign T76 = ~ T77;
  assign T77 = T78[9];
  assign T78 = T79 - 13'h310;
  assign T79 = $signed(io_in_19) * $signed(3'h2);
  assign io_out_20 = T80;
  assign T80 = ~ T81;
  assign T81 = T82[9];
  assign T82 = T83 - 13'h310;
  assign T83 = $signed(io_in_20) * $signed(3'h2);
  assign io_out_21 = T84;
  assign T84 = ~ T85;
  assign T85 = T86[9];
  assign T86 = T87 - 13'h310;
  assign T87 = $signed(io_in_21) * $signed(3'h2);
  assign io_out_22 = T88;
  assign T88 = ~ T89;
  assign T89 = T90[9];
  assign T90 = T91 - 13'h310;
  assign T91 = $signed(io_in_22) * $signed(3'h2);
  assign io_out_23 = T92;
  assign T92 = ~ T93;
  assign T93 = T94[9];
  assign T94 = T95 - 13'h310;
  assign T95 = $signed(io_in_23) * $signed(3'h2);
  assign io_out_24 = T96;
  assign T96 = ~ T97;
  assign T97 = T98[9];
  assign T98 = T99 - 13'h310;
  assign T99 = $signed(io_in_24) * $signed(3'h2);
  assign io_out_25 = T100;
  assign T100 = ~ T101;
  assign T101 = T102[9];
  assign T102 = T103 - 13'h310;
  assign T103 = $signed(io_in_25) * $signed(3'h2);
  assign io_out_26 = T104;
  assign T104 = ~ T105;
  assign T105 = T106[9];
  assign T106 = T107 - 13'h310;
  assign T107 = $signed(io_in_26) * $signed(3'h2);
  assign io_out_27 = T108;
  assign T108 = ~ T109;
  assign T109 = T110[9];
  assign T110 = T111 - 13'h310;
  assign T111 = $signed(io_in_27) * $signed(3'h2);
  assign io_out_28 = T112;
  assign T112 = ~ T113;
  assign T113 = T114[9];
  assign T114 = T115 - 13'h310;
  assign T115 = $signed(io_in_28) * $signed(3'h2);
  assign io_out_29 = T116;
  assign T116 = ~ T117;
  assign T117 = T118[9];
  assign T118 = T119 - 13'h310;
  assign T119 = $signed(io_in_29) * $signed(3'h2);
  assign io_out_30 = T120;
  assign T120 = ~ T121;
  assign T121 = T122[9];
  assign T122 = T123 - 13'h310;
  assign T123 = $signed(io_in_30) * $signed(3'h2);
  assign io_out_31 = T124;
  assign T124 = ~ T125;
  assign T125 = T126[9];
  assign T126 = T127 - 13'h310;
  assign T127 = $signed(io_in_31) * $signed(3'h2);
endmodule

module MemoryUnit_0(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T5;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T6;
  reg  restartRegs_0;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (addr)
    0: T0 = 32'h13077655;
    1: T0 = 32'h7ff288b;
    2: T0 = 32'h5d200573;
    3: T0 = 32'hbb4149ed;
    4: T0 = 32'h62591000;
    5: T0 = 32'hf3ff0419;
    6: T0 = 32'h39e07440;
    7: T0 = 32'h53ff1413;
    8: T0 = 32'hc63a61d8;
    9: T0 = 32'hc6bdfffd;
    10: T0 = 32'hc1aae042;
    11: T0 = 32'h12e06010;
    12: T0 = 32'hf870ad6;
    13: T0 = 32'h10d84000;
    14: T0 = 32'hc0180073;
    15: T0 = 32'h4bc5800;
    16: T0 = 32'hf800f00a;
    17: T0 = 32'he785ff;
    18: T0 = 32'hfc80ffff;
    19: T0 = 32'h1fff93;
    20: T0 = 32'hfffebfff;
    21: T0 = 32'h33ffffff;
    22: T0 = 32'hfdf8e7ff;
    23: T0 = 32'hc21fc1ff;
    24: T0 = 32'hffcffaef;
    25: T0 = 32'h1cb5e00b;
    26: T0 = 32'ha7f81ff7;
    27: T0 = 32'h80f68602;
    28: T0 = 32'hf7ff1fbe;
    29: T0 = 32'he00ccc00;
    30: T0 = 32'h37ff03e4;
    31: T0 = 32'hf800e4d0;
    32: T0 = 32'h7b3f003e;
    33: T0 = 32'h1f00f826;
    34: T0 = 32'h3b71b004;
    35: T0 = 32'h5bf0e4c7;
    36: T0 = 32'h7f76601;
    37: T0 = 32'hd16eff2e;
    38: T0 = 32'he2136d2b;
    39: T0 = 32'h79f1ffbe;
    40: T0 = 32'hde063dd2;
    41: T0 = 32'h670207ff;
    42: T0 = 32'h5fc0ac38;
    43: T0 = 32'hd932d7e;
    44: T0 = 32'h27be8016;
    45: T0 = 32'he55b3b27;
    46: T0 = 32'hf237abe3;
    47: T0 = 32'h5feee70f;
    48: T0 = 32'h22898807;
    49: T0 = 32'h2e4cd646;
    50: T0 = 32'h26b52e7d;
    51: T0 = 32'h54a35553;
    52: T0 = 32'h6a0323b6;
    53: T0 = 32'h2caa41e4;
    54: T0 = 32'hb92d0ad8;
    55: T0 = 32'hca876ae9;
    56: T0 = 32'h56804200;
    57: T0 = 32'h403158f0;
    58: T0 = 32'h94d80015;
    59: T0 = 32'he700da1e;
    60: T0 = 32'h11bfff7f;
    61: T0 = 32'he03cfeaf;
    62: T0 = 32'he1037fff;
    63: T0 = 32'hdf03fbec;
    64: T0 = 32'h3e0f79ff;
    65: T0 = 32'he3f8fbfc;
    66: T0 = 32'h83e0110f;
    67: T0 = 32'h5b85f3a;
    68: T0 = 32'hc43ff0b8;
    69: T0 = 32'he09d8f13;
    70: T0 = 32'h80c33fc7;
    71: T0 = 32'h3f037fc3;
    72: T0 = 32'h4ac401fe;
    73: T0 = 32'h3c8fbc6;
    74: T0 = 32'h71fca0f;
    75: T0 = 32'hd03cff60;
    76: T0 = 32'he0af09f0;
    77: T0 = 32'hfdc317f2;
    78: T0 = 32'h1f83204e;
    79: T0 = 32'h777eebb4;
    80: T0 = 32'he1fc0684;
    81: T0 = 32'hc6831000;
    82: T0 = 32'h199f0014;
    83: T0 = 32'hfc18c200;
    84: T0 = 32'h80090004;
    85: T0 = 32'h1fc4cc28;
    86: T0 = 32'h100000;
    87: T0 = 32'h1fc2382;
    88: T0 = 32'hd0a163f0;
    89: T0 = 32'h1ffe9c;
    90: T0 = 32'h9002abff;
    91: T0 = 32'h200bffe8;
    92: T0 = 32'h7c33295f;
    93: T0 = 32'h58c1ffff;
    94: T0 = 32'h80437a64;
    95: T0 = 32'h198eda32;
    96: T0 = 32'h7fb06c05;
    97: T0 = 32'h81736b91;
    98: T0 = 32'h43b7326c;
    99: T0 = 32'h7777058b;
    100: T0 = 32'h9f85a4e5;
    101: T0 = 32'h8e85eb3c;
    102: T0 = 32'h368ec03a;
    103: T0 = 32'h40e14ed2;
    104: T0 = 32'he5ca1f80;
    105: T0 = 32'ha8011f03;
    106: T0 = 32'h5fe11bfe;
    107: T0 = 32'hcf82fdf1;
    108: T0 = 32'h3eba6ff;
    109: T0 = 32'h6b60ffd7;
    110: T0 = 32'hcd7c37;
    111: T0 = 32'hd8f66080;
    112: T0 = 32'hd0270bfc;
    113: T0 = 32'hff820000;
    114: T0 = 32'h37fb01fe;
    115: T0 = 32'hfc70f100;
    116: T0 = 32'h9ff001f;
    117: T0 = 32'hb3c0ff8e;
    118: T0 = 32'hd7e0b1;
    119: T0 = 32'hf0101d38;
    120: T0 = 32'h971e;
    121: T0 = 32'hf600f0c2;
    122: T0 = 32'h3453;
    123: T0 = 32'hae0df04;
    124: T0 = 32'h60387a;
    125: T0 = 32'he03efbfc;
    126: T0 = 32'he017e106;
    127: T0 = 32'hffe19e3f;
    128: T0 = 32'h4b20ff03;
    129: T0 = 32'hffe6278;
    130: T0 = 32'he4f581f0;
    131: T0 = 32'ha07f0210;
    132: T0 = 32'hbec3181f;
    133: T0 = 32'h7a070036;
    134: T0 = 32'h39e852c0;
    135: T0 = 32'hbb001060;
    136: T0 = 32'hc0ff069f;
    137: T0 = 32'h7294f407;
    138: T0 = 32'h5c07a089;
    139: T0 = 32'h1e47f04;
    140: T0 = 32'h200000c3;
    141: T0 = 32'h24317c;
    142: T0 = 32'hb400001e;
    143: T0 = 32'h700512ae;
    144: T0 = 32'hdb8c8003;
    145: T0 = 32'h425336be;
    146: T0 = 32'ha9acccaf;
    147: T0 = 32'he6918de1;
    148: T0 = 32'h778180ef;
    149: T0 = 32'h3fa21276;
    150: T0 = 32'h2a7c4b62;
    151: T0 = 32'he01b3b2f;
    152: T0 = 32'hb640e5a5;
    153: T0 = 32'h342e007f;
    154: T0 = 32'hcd01ffc7;
    155: T0 = 32'hfa8fa000;
    156: T0 = 32'ha5410342;
    157: T0 = 32'hfffb19c0;
    158: T0 = 32'hfea07000;
    159: T0 = 32'hffff0057;
    160: T0 = 32'hffe7e000;
    161: T0 = 32'h7fff8007;
    162: T0 = 32'hfff77600;
    163: T0 = 32'hc7ff3c01;
    164: T0 = 32'hffff9d10;
    165: T0 = 32'he3ff85c0;
    166: T0 = 32'hfe1f06ed;
    167: T0 = 32'h6177e2e;
    168: T0 = 32'h9c00e02f;
    169: T0 = 32'h358f8;
    170: T0 = 32'h70f8e700;
    171: T0 = 32'hd0008abf;
    172: T0 = 32'h2a1f0f9;
    173: T0 = 32'h3c804527;
    174: T0 = 32'h38679c6;
    175: T0 = 32'h4bc0603e;
    176: T0 = 32'h102887e5;
    177: T0 = 32'h18aff0df;
    178: T0 = 32'hf107743e;
    179: T0 = 32'he484e7ff;
    180: T0 = 32'h908ff4f;
    181: T0 = 32'h1f13ffff;
    182: T0 = 32'h4130fffc;
    183: T0 = 32'he7ee3b37;
    184: T0 = 32'haf780fff;
    185: T0 = 32'hfffef430;
    186: T0 = 32'hd86f0006;
    187: T0 = 32'h7fff065e;
    188: T0 = 32'hf86ad000;
    189: T0 = 32'h9d3f0009;
    190: T0 = 32'hfc46a480;
    191: T0 = 32'ha51f4000;
    192: T0 = 32'h7fa0d318;
    193: T0 = 32'hfed6443;
    194: T0 = 32'ha341cd4f;
    195: T0 = 32'h52b753af;
    196: T0 = 32'hbd51a0d4;
    197: T0 = 32'h5e2a7778;
    198: T0 = 32'h642017ed;
    199: T0 = 32'hec52c59c;
    200: T0 = 32'h697323c9;
    201: T0 = 32'h25010011;
    202: T0 = 32'h111bd8b8;
    203: T0 = 32'h5f00c141;
    204: T0 = 32'h156477b;
    205: T0 = 32'h3d4078fe;
    206: T0 = 32'h80f7d87b;
    207: T0 = 32'hfedff70f;
    208: T0 = 32'he0ffe07c;
    209: T0 = 32'hfd6b27f1;
    210: T0 = 32'h201f9f0d;
    211: T0 = 32'hffb40c3f;
    212: T0 = 32'hed0178fc;
    213: T0 = 32'h7ff12280;
    214: T0 = 32'hc8d80387;
    215: T0 = 32'h87ff0022;
    216: T0 = 32'h5bfa038;
    217: T0 = 32'h40700000;
    218: T0 = 32'h653303;
    219: T0 = 32'hff823000;
    220: T0 = 32'h2050a00;
    221: T0 = 32'he7e8300;
    222: T0 = 32'hf09fc049;
    223: T0 = 32'hfe770030;
    224: T0 = 32'h1f01ff02;
    225: T0 = 32'h3ec121e1;
    226: T0 = 32'hb7f81ffe;
    227: T0 = 32'hc3aef67f;
    228: T0 = 32'h47ffc07f;
    229: T0 = 32'hff00efb7;
    230: T0 = 32'h2bca07;
    231: T0 = 32'h7ff03f1f;
    232: T0 = 32'h8004fbbc;
    233: T0 = 32'h157f81d7;
    234: T0 = 32'h9400fc5f;
    235: T0 = 32'h6c95f861;
    236: T0 = 32'h80300629;
    237: T0 = 32'hff7c0000;
    238: T0 = 32'h100700ec;
    239: T0 = 32'hffc4fa00;
    240: T0 = 32'h97dc0eaf;
    241: T0 = 32'hffe1a236;
    242: T0 = 32'h3e2b61c7;
    243: T0 = 32'h3ffc797e;
    244: T0 = 32'h9fc3ea59;
    245: T0 = 32'h2c9b6f80;
    246: T0 = 32'hf5c20ef5;
    247: T0 = 32'h368867f5;
    248: T0 = 32'hb155202a;
    249: T0 = 32'ha3930f9;
    250: T0 = 32'hc352f61d;
    251: T0 = 32'hd713f7f7;
    252: T0 = 32'h90071fce;
    253: T0 = 32'h7fa697fc;
    254: T0 = 32'h3c00007c;
    255: T0 = 32'h786ffd8;
    256: T0 = 32'hfe400007;
    257: T0 = 32'h7e01f3e;
    258: T0 = 32'h7ad7000;
    259: T0 = 32'h6bff00fe;
    260: T0 = 32'hf0737a6e;
    261: T0 = 32'hd3fffc01;
    262: T0 = 32'hff071b2f;
    263: T0 = 32'h73ff7ff0;
    264: T0 = 32'hdff0c05f;
    265: T0 = 32'h78f201f;
    266: T0 = 32'hffee3f08;
    267: T0 = 32'he7f67410;
    268: T0 = 32'hf21cf3fd;
    269: T0 = 32'h477ff833;
    270: T0 = 32'hf7a1bf3f;
    271: T0 = 32'hc67efab;
    272: T0 = 32'h3fe49ff9;
    273: T0 = 32'he0c28fea;
    274: T0 = 32'hfcefbf;
    275: T0 = 32'hfd44f86d;
    276: T0 = 32'h700f4c6f;
    277: T0 = 32'h7ab4efdc;
    278: T0 = 32'hff808039;
    279: T0 = 32'h7f5afff;
    280: T0 = 32'h7ff8c01b;
    281: T0 = 32'h72e6af;
    282: T0 = 32'he7df0301;
    283: T0 = 32'hf0037ca0;
    284: T0 = 32'h7880010;
    285: T0 = 32'h7e20e81c;
    286: T0 = 32'h720f4401;
    287: T0 = 32'h9be10e08;
    288: T0 = 32'h621f4d20;
    289: T0 = 32'h37dc01e0;
    290: T0 = 32'h16b0edd4;
    291: T0 = 32'h34cbe1ff;
    292: T0 = 32'h8c8bb6;
    293: T0 = 32'h3b39a52a;
    294: T0 = 32'hda494eda;
    295: T0 = 32'hb48e9bb8;
    296: T0 = 32'ha0ca7727;
    297: T0 = 32'hd2a0ca79;
    298: T0 = 32'h83732ff7;
    299: T0 = 32'h7f1afda0;
    300: T0 = 32'hd433fff;
    301: T0 = 32'h4ffffffc;
    302: T0 = 32'h20d42bff;
    303: T0 = 32'h30fcffff;
    304: T0 = 32'hf85bfa9f;
    305: T0 = 32'h95f3fff;
    306: T0 = 32'hffc1fe94;
    307: T0 = 32'h1c540ff;
    308: T0 = 32'h8dfcffcf;
    309: T0 = 32'h250e01;
    310: T0 = 32'hc0050010;
    311: T0 = 32'h80000e48;
    312: T0 = 32'h7d011000;
    313: T0 = 32'h3c0478;
    314: T0 = 32'hfee8d1c4;
    315: T0 = 32'h9fe7600d;
    316: T0 = 32'hfffe13ff;
    317: T0 = 32'h99ffde00;
    318: T0 = 32'hfffe291f;
    319: T0 = 32'hfabfece0;
    320: T0 = 32'hffff0187;
    321: T0 = 32'hffc14f4e;
    322: T0 = 32'h9ffc7c57;
    323: T0 = 32'h81ffe810;
    324: T0 = 32'h19ef0041;
    325: T0 = 32'hf00700c4;
    326: T0 = 32'h3baf7f3d;
    327: T0 = 32'hff00fab8;
    328: T0 = 32'h410fff;
    329: T0 = 32'h5ff0ffe4;
    330: T0 = 32'h601d17f;
    331: T0 = 32'hb56f7fff;
    332: T0 = 32'hf338fa07;
    333: T0 = 32'h310d1fff;
    334: T0 = 32'hdd607f3a;
    335: T0 = 32'h804f03fc;
    336: T0 = 32'h2eaf5e5;
    337: T0 = 32'hc6b0037e;
    338: T0 = 32'hb2ff3dfe;
    339: T0 = 32'hf82c27bc;
    340: T0 = 32'hdf9b0815;
    341: T0 = 32'h2771fe82;
    342: T0 = 32'he6844c70;
    343: T0 = 32'h12a6c978;
    344: T0 = 32'h6bc7e688;
    345: T0 = 32'h8c1e9f1d;
    346: T0 = 32'hbff06565;
    347: T0 = 32'h6657c283;
    348: T0 = 32'h7f7c26ba;
    349: T0 = 32'h7d135e2;
    350: T0 = 32'hbffe06d6;
    351: T0 = 32'h2caafe;
    352: T0 = 32'h2ffafc7e;
    353: T0 = 32'h810673af;
    354: T0 = 32'h9fc3fe0;
    355: T0 = 32'h9f80071a;
    356: T0 = 32'h2e681ff;
    357: T0 = 32'h47fcf07a;
    358: T0 = 32'hf03dbc03;
    359: T0 = 32'ha91f0f06;
    360: T0 = 32'h7c05340;
    361: T0 = 32'h194000e0;
    362: T0 = 32'h1e0930;
    363: T0 = 32'he074018e;
    364: T0 = 32'h2e095;
    365: T0 = 32'h3e06ca1f;
    366: T0 = 32'he4007e00;
    367: T0 = 32'hc7e01841;
    368: T0 = 32'h6010d70;
    369: T0 = 32'h383ec7ec;
    370: T0 = 32'he0f4bbf2;
    371: T0 = 32'h3c1be1d;
    372: T0 = 32'h1e062bff;
    373: T0 = 32'h3c1cf8f8;
    374: T0 = 32'hf0c19c48;
    375: T0 = 32'h2041b387;
    376: T0 = 32'hf8c396a;
    377: T0 = 32'h8f089b18;
    378: T0 = 32'hc0f5c398;
    379: T0 = 32'h7cd1aaed;
    380: T0 = 32'hc01cf439;
    381: T0 = 32'h6fd0c698;
    382: T0 = 32'hd88ea17;
    383: T0 = 32'h3f1fe09;
    384: T0 = 32'h78316bc0;
    385: T0 = 32'ha3800fd9;
    386: T0 = 32'hf41df03c;
    387: T0 = 32'hac06fffb;
    388: T0 = 32'h3fffcc6e;
    389: T0 = 32'h3df4adff;
    390: T0 = 32'h62fd3e81;
    391: T0 = 32'h3fecd1e5;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T5 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T6 = reset ? 1'h0 : restartRegs_0;
  assign T7 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_1(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T5;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T6;
  reg  restartRegs_0;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (addr)
    0: T0 = 32'ha396095f;
    1: T0 = 32'hf1bc1aa8;
    2: T0 = 32'hc05df887;
    3: T0 = 32'h34b4c215;
    4: T0 = 32'h9d079df7;
    5: T0 = 32'hc9ffed9d;
    6: T0 = 32'hffd2b3ef;
    7: T0 = 32'h200b210b;
    8: T0 = 32'h5fc969f3;
    9: T0 = 32'h99c4a357;
    10: T0 = 32'hffffe03f;
    11: T0 = 32'hf2f2ffff;
    12: T0 = 32'he07ff153;
    13: T0 = 32'hffe50fff;
    14: T0 = 32'h4801ffde;
    15: T0 = 32'h7f9f03f;
    16: T0 = 32'ha200d33e;
    17: T0 = 32'hf03f6202;
    18: T0 = 32'hfe8fedf7;
    19: T0 = 32'h7f80e720;
    20: T0 = 32'h3fdcf7f;
    21: T0 = 32'hfff1f6f0;
    22: T0 = 32'h1c349bff;
    23: T0 = 32'h8bebfe1b;
    24: T0 = 32'h1e7318f;
    25: T0 = 32'hf1ff3ee0;
    26: T0 = 32'hf80f01cf;
    27: T0 = 32'h3a13484c;
    28: T0 = 32'h7ff84016;
    29: T0 = 32'h80b8e800;
    30: T0 = 32'h7fff8201;
    31: T0 = 32'hfc0c0881;
    32: T0 = 32'hea4f0000;
    33: T0 = 32'h1fc0014c;
    34: T0 = 32'hdc8a000;
    35: T0 = 32'hfe0008;
    36: T0 = 32'hfcde5400;
    37: T0 = 32'hc60700b8;
    38: T0 = 32'h1d146e0;
    39: T0 = 32'h88003ff2;
    40: T0 = 32'h3e4ce;
    41: T0 = 32'h9162f3ff;
    42: T0 = 32'h3bbeffbd;
    43: T0 = 32'h7ee825ff;
    44: T0 = 32'hfa3efffe;
    45: T0 = 32'h800636a7;
    46: T0 = 32'h2cb78087;
    47: T0 = 32'h6081f9bb;
    48: T0 = 32'hb0a666b6;
    49: T0 = 32'hd4267f06;
    50: T0 = 32'h52463ceb;
    51: T0 = 32'h1b25f8aa;
    52: T0 = 32'haaf879a4;
    53: T0 = 32'hcdc0f880;
    54: T0 = 32'h77d24354;
    55: T0 = 32'h51d73c07;
    56: T0 = 32'h8ffa7f62;
    57: T0 = 32'hb600f00;
    58: T0 = 32'hb4b81dae;
    59: T0 = 32'h48fe7ce0;
    60: T0 = 32'hfc8e017f;
    61: T0 = 32'h800fc746;
    62: T0 = 32'h3f98103e;
    63: T0 = 32'h3d00e0fc;
    64: T0 = 32'hba2007;
    65: T0 = 32'hc2007e06;
    66: T0 = 32'h80003a60;
    67: T0 = 32'h3e203e0;
    68: T0 = 32'h378001d4;
    69: T0 = 32'h80d01f;
    70: T0 = 32'h801cfa0f;
    71: T0 = 32'hf0008701;
    72: T0 = 32'hc0011f81;
    73: T0 = 32'h1fd00c70;
    74: T0 = 32'hfbb980e6;
    75: T0 = 32'hd9ff1484;
    76: T0 = 32'hffd0761f;
    77: T0 = 32'hafff60c3;
    78: T0 = 32'hfffd07f8;
    79: T0 = 32'hd97ec600;
    80: T0 = 32'hdfff053f;
    81: T0 = 32'h3f3ffd40;
    82: T0 = 32'h65fa0005;
    83: T0 = 32'he1761ff0;
    84: T0 = 32'h607f0a00;
    85: T0 = 32'h500d17bc;
    86: T0 = 32'h1e07c840;
    87: T0 = 32'h1bb;
    88: T0 = 32'h2ef03706;
    89: T0 = 32'h80f046;
    90: T0 = 32'h47da34c1;
    91: T0 = 32'ha0000f09;
    92: T0 = 32'h3f6cc7b4;
    93: T0 = 32'h622046e2;
    94: T0 = 32'h1429da1;
    95: T0 = 32'h23609b81;
    96: T0 = 32'h800079e9;
    97: T0 = 32'h16c7089c;
    98: T0 = 32'h2f1f5a42;
    99: T0 = 32'h88fc2627;
    100: T0 = 32'hb07b4c6f;
    101: T0 = 32'he6184c49;
    102: T0 = 32'h874769e4;
    103: T0 = 32'hec4750fe;
    104: T0 = 32'hf0ed5e00;
    105: T0 = 32'hb68f0035;
    106: T0 = 32'hff4ac5ff;
    107: T0 = 32'h84d7fc2d;
    108: T0 = 32'hfefdf43d;
    109: T0 = 32'h7b79ffff;
    110: T0 = 32'hd17fff37;
    111: T0 = 32'hfeed7fff;
    112: T0 = 32'h77ffffe2;
    113: T0 = 32'hfb63d3ff;
    114: T0 = 32'h4a5fc3bf;
    115: T0 = 32'h7c006a9f;
    116: T0 = 32'h151783f;
    117: T0 = 32'hf6f3;
    118: T0 = 32'h2e57053;
    119: T0 = 32'hd8409feb;
    120: T0 = 32'h47bd707;
    121: T0 = 32'hd1078ff;
    122: T0 = 32'hc073bf40;
    123: T0 = 32'h94014e03;
    124: T0 = 32'h1f24;
    125: T0 = 32'h17046f0;
    126: T0 = 32'hc18097a3;
    127: T0 = 32'h9a073;
    128: T0 = 32'h104889a8;
    129: T0 = 32'h10280;
    130: T0 = 32'h3a401800;
    131: T0 = 32'h6000068;
    132: T0 = 32'h75a2200;
    133: T0 = 32'hb7fc0007;
    134: T0 = 32'hffee7c02;
    135: T0 = 32'h90dfff00;
    136: T0 = 32'hffff847d;
    137: T0 = 32'he9177fff;
    138: T0 = 32'hbeffffa9;
    139: T0 = 32'hfc81afff;
    140: T0 = 32'he61fffc;
    141: T0 = 32'hfbf570af;
    142: T0 = 32'h58c7bff9;
    143: T0 = 32'h3fff30d8;
    144: T0 = 32'hc2c7ceb1;
    145: T0 = 32'h42fc4379;
    146: T0 = 32'hcd33d133;
    147: T0 = 32'h37054eec;
    148: T0 = 32'h130fedd7;
    149: T0 = 32'h82677f94;
    150: T0 = 32'h243e6c4d;
    151: T0 = 32'h319a01ff;
    152: T0 = 32'h2b01eb52;
    153: T0 = 32'h1465a03f;
    154: T0 = 32'h41fcfd93;
    155: T0 = 32'h881c7003;
    156: T0 = 32'h14df0fcd;
    157: T0 = 32'hf83c0cfc;
    158: T0 = 32'hb20a6c3f;
    159: T0 = 32'h2fe2f8c4;
    160: T0 = 32'h80d007c1;
    161: T0 = 32'h86ff1f9f;
    162: T0 = 32'hf02edc06;
    163: T0 = 32'hfb5fe1f2;
    164: T0 = 32'h9e41e4ce;
    165: T0 = 32'hafdbb1f;
    166: T0 = 32'hf0e5f4a8;
    167: T0 = 32'h1827bef1;
    168: T0 = 32'hfc0e0f90;
    169: T0 = 32'hf380bdd7;
    170: T0 = 32'hb7d020fe;
    171: T0 = 32'hf30ecbf;
    172: T0 = 32'h3f70ed83;
    173: T0 = 32'h4780e07;
    174: T0 = 32'hc3871e44;
    175: T0 = 32'h780360ff;
    176: T0 = 32'h3c7501d0;
    177: T0 = 32'h8cc08307;
    178: T0 = 32'h81e63191;
    179: T0 = 32'h6462478;
    180: T0 = 32'h601fc3e1;
    181: T0 = 32'hf1829663;
    182: T0 = 32'h8f417c16;
    183: T0 = 32'h4fdc3b4e;
    184: T0 = 32'hd87f07c3;
    185: T0 = 32'hffbf3074;
    186: T0 = 32'h7a6343e8;
    187: T0 = 32'haff887a9;
    188: T0 = 32'h9ff1b2bf;
    189: T0 = 32'h9afbf051;
    190: T0 = 32'hf538a600;
    191: T0 = 32'h2a05f8fd;
    192: T0 = 32'hfe27a72f;
    193: T0 = 32'hda1c3b77;
    194: T0 = 32'hfed6a37a;
    195: T0 = 32'h786bf6d;
    196: T0 = 32'h1e13649c;
    197: T0 = 32'hc43012d4;
    198: T0 = 32'hbc58dde5;
    199: T0 = 32'h97942440;
    200: T0 = 32'hd05d9196;
    201: T0 = 32'hb318d1b9;
    202: T0 = 32'h488f8977;
    203: T0 = 32'hfbe41df0;
    204: T0 = 32'h2fcbc098;
    205: T0 = 32'hb449001e;
    206: T0 = 32'h3ffe895c;
    207: T0 = 32'hf2400000;
    208: T0 = 32'h2c0100dc;
    209: T0 = 32'h2fe7343e;
    210: T0 = 32'h7fe0c81b;
    211: T0 = 32'h95e812;
    212: T0 = 32'hbbff0000;
    213: T0 = 32'hfe0008e0;
    214: T0 = 32'h148f0000;
    215: T0 = 32'hf8781067;
    216: T0 = 32'hf8487808;
    217: T0 = 32'h9f03e08d;
    218: T0 = 32'h1fe2e7e1;
    219: T0 = 32'h39e0ffff;
    220: T0 = 32'hc1fff03f;
    221: T0 = 32'hf42effff;
    222: T0 = 32'hdbffffb7;
    223: T0 = 32'hff3bdfff;
    224: T0 = 32'h4c0ffffd;
    225: T0 = 32'h7ff5c637;
    226: T0 = 32'he0c17fff;
    227: T0 = 32'h7bf8f5d8;
    228: T0 = 32'h1850aff;
    229: T0 = 32'h7f8fff8c;
    230: T0 = 32'hb5c107;
    231: T0 = 32'h2ff85c02;
    232: T0 = 32'he0022601;
    233: T0 = 32'hdcf60000;
    234: T0 = 32'h6f801de0;
    235: T0 = 32'hf004000;
    236: T0 = 32'h137c0068;
    237: T0 = 32'he36ae580;
    238: T0 = 32'ha15f00bb;
    239: T0 = 32'h7fee5a7e;
    240: T0 = 32'h12a1ffc2;
    241: T0 = 32'h1f18bdf;
    242: T0 = 32'hf260a9f8;
    243: T0 = 32'h201ec937;
    244: T0 = 32'h8d2c0da6;
    245: T0 = 32'h9c572bb0;
    246: T0 = 32'h2b342296;
    247: T0 = 32'h56c6ffb9;
    248: T0 = 32'h5472d696;
    249: T0 = 32'h5c3f691d;
    250: T0 = 32'hffe0dc90;
    251: T0 = 32'hc7ccd2f7;
    252: T0 = 32'h3ffff87e;
    253: T0 = 32'hfeac8b0f;
    254: T0 = 32'h5fff8b2;
    255: T0 = 32'hfffdf4e0;
    256: T0 = 32'hb5c33f07;
    257: T0 = 32'h1b0b60;
    258: T0 = 32'h3f20a3e0;
    259: T0 = 32'h100;
    260: T0 = 32'h11f225fe;
    261: T0 = 32'hf4008010;
    262: T0 = 32'h17ff1e7f;
    263: T0 = 32'heec0f010;
    264: T0 = 32'he7fff05b;
    265: T0 = 32'hfb307f03;
    266: T0 = 32'h3fe73f02;
    267: T0 = 32'h1f0564f8;
    268: T0 = 32'hbffec1ff;
    269: T0 = 32'h2000c10f;
    270: T0 = 32'h71c3e9f;
    271: T0 = 32'he0007ca4;
    272: T0 = 32'h757e9;
    273: T0 = 32'hff8093f4;
    274: T0 = 32'h401c1ff;
    275: T0 = 32'h4279f81e;
    276: T0 = 32'hb0f0f83a;
    277: T0 = 32'ha03ec3c1;
    278: T0 = 32'hfb1f1eb4;
    279: T0 = 32'hff9d8e9e;
    280: T0 = 32'h9feff3f2;
    281: T0 = 32'hfff938fc;
    282: T0 = 32'h73676f2b;
    283: T0 = 32'hffff98a4;
    284: T0 = 32'hf3f0787f;
    285: T0 = 32'h9ff440;
    286: T0 = 32'hee3a10d3;
    287: T0 = 32'h2af9f4b;
    288: T0 = 32'h7fa86417;
    289: T0 = 32'h365341fd;
    290: T0 = 32'hfdfec529;
    291: T0 = 32'hbc83080c;
    292: T0 = 32'h4f7bab45;
    293: T0 = 32'h1071cb2b;
    294: T0 = 32'h54db3214;
    295: T0 = 32'h2d045219;
    296: T0 = 32'hf41f31e;
    297: T0 = 32'h66d095bf;
    298: T0 = 32'hccfb7f9f;
    299: T0 = 32'h1fb450df;
    300: T0 = 32'ha24e9000;
    301: T0 = 32'hecff4c5e;
    302: T0 = 32'hff399900;
    303: T0 = 32'ha3372326;
    304: T0 = 32'hd3fecdd6;
    305: T0 = 32'hf7d2bff0;
    306: T0 = 32'h3be5f;
    307: T0 = 32'hfa16bfe;
    308: T0 = 32'h2800e172;
    309: T0 = 32'h3f0407;
    310: T0 = 32'h7ba0087a;
    311: T0 = 32'hf0019280;
    312: T0 = 32'h9790003;
    313: T0 = 32'h7fe07fa8;
    314: T0 = 32'hc0ef8008;
    315: T0 = 32'he303ffe1;
    316: T0 = 32'h3f095034;
    317: T0 = 32'h98006ffc;
    318: T0 = 32'h1fcc6c0;
    319: T0 = 32'hec7c83ff;
    320: T0 = 32'hf01ff071;
    321: T0 = 32'hffcdde1f;
    322: T0 = 32'hbfe8f807;
    323: T0 = 32'h87fc79a3;
    324: T0 = 32'hcfff7000;
    325: T0 = 32'h786f07c6;
    326: T0 = 32'h8dffdf00;
    327: T0 = 32'h6f8400dc;
    328: T0 = 32'hf03ce5f0;
    329: T0 = 32'h917f0038;
    330: T0 = 32'hfe0cd36f;
    331: T0 = 32'h422de65f;
    332: T0 = 32'h7180f813;
    333: T0 = 32'heb403e1f;
    334: T0 = 32'hc9cff8c;
    335: T0 = 32'hff2b79e7;
    336: T0 = 32'hb5021ffe;
    337: T0 = 32'hf97a473e;
    338: T0 = 32'h4a39d7fe;
    339: T0 = 32'h7d5d7;
    340: T0 = 32'hcd02407f;
    341: T0 = 32'h6806ed6d;
    342: T0 = 32'hc864ded;
    343: T0 = 32'h6c85da6a;
    344: T0 = 32'hce32ec4;
    345: T0 = 32'h4c3137bc;
    346: T0 = 32'h60a0c1b0;
    347: T0 = 32'h22f69340;
    348: T0 = 32'hbf631f0a;
    349: T0 = 32'habc63068;
    350: T0 = 32'h303c6467;
    351: T0 = 32'heb46eedc;
    352: T0 = 32'h7301fff9;
    353: T0 = 32'hf39bd5f;
    354: T0 = 32'hc9c8f81f;
    355: T0 = 32'hc03f2e3f;
    356: T0 = 32'hff4b7fc0;
    357: T0 = 32'hcf0003bd;
    358: T0 = 32'hfff77fc;
    359: T0 = 32'h6440e0fe;
    360: T0 = 32'h203fec3f;
    361: T0 = 32'hf5837e1f;
    362: T0 = 32'hb0ffecf;
    363: T0 = 32'hffc05471;
    364: T0 = 32'hdc7108e5;
    365: T0 = 32'hff5ee1f;
    366: T0 = 32'hb3e7fb81;
    367: T0 = 32'hb0e70a61;
    368: T0 = 32'hff5f1ef8;
    369: T0 = 32'hef01004c;
    370: T0 = 32'h1c2f805f;
    371: T0 = 32'haff8e010;
    372: T0 = 32'he0f8d003;
    373: T0 = 32'hd0d11a00;
    374: T0 = 32'h7f01f950;
    375: T0 = 32'h14308830;
    376: T0 = 32'h678ffff;
    377: T0 = 32'h808b7821;
    378: T0 = 32'h11670ff8;
    379: T0 = 32'hf83b23ef;
    380: T0 = 32'h318280ff;
    381: T0 = 32'h2781eaef;
    382: T0 = 32'h1e387c6f;
    383: T0 = 32'h1807e3e;
    384: T0 = 32'h2e75dbde;
    385: T0 = 32'he67c43fb;
    386: T0 = 32'h20ebc191;
    387: T0 = 32'h996f001e;
    388: T0 = 32'hcffce4b8;
    389: T0 = 32'h5d848082;
    390: T0 = 32'hd8394f25;
    391: T0 = 32'h3e3be34;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T5 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T6 = reset ? 1'h0 : restartRegs_0;
  assign T7 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_2(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T5;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T6;
  reg  restartRegs_0;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (addr)
    0: T0 = 32'h1edeba33;
    1: T0 = 32'h480dfff;
    2: T0 = 32'h9fa5f9fb;
    3: T0 = 32'h74260554;
    4: T0 = 32'h8e201189;
    5: T0 = 32'hf8d3a052;
    6: T0 = 32'h266c000;
    7: T0 = 32'hfee0f81d;
    8: T0 = 32'h60f083;
    9: T0 = 32'hb840ffe8;
    10: T0 = 32'h1e13f;
    11: T0 = 32'h10e0f007;
    12: T0 = 32'h90f37;
    13: T0 = 32'hfd487e80;
    14: T0 = 32'h703f000f;
    15: T0 = 32'hffda17fc;
    16: T0 = 32'h3ffff000;
    17: T0 = 32'hfffe06fe;
    18: T0 = 32'h7dff4f80;
    19: T0 = 32'hffff0054;
    20: T0 = 32'he7bfc43c;
    21: T0 = 32'h3efff800;
    22: T0 = 32'hc0c14238;
    23: T0 = 32'hce00c7fb;
    24: T0 = 32'h1f8c3;
    25: T0 = 32'h2a03e7f;
    26: T0 = 32'hf1107e3b;
    27: T0 = 32'hf15932cf;
    28: T0 = 32'h6a09f3fd;
    29: T0 = 32'h19d287bf;
    30: T0 = 32'h78407f0f;
    31: T0 = 32'h7a26766a;
    32: T0 = 32'hfbcc00e0;
    33: T0 = 32'hce6907e4;
    34: T0 = 32'h39ff2000;
    35: T0 = 32'hef80007c;
    36: T0 = 32'hf440;
    37: T0 = 32'hfb201001;
    38: T0 = 32'h1740;
    39: T0 = 32'h5f8cc00;
    40: T0 = 32'he570;
    41: T0 = 32'hb225fff;
    42: T0 = 32'h8012;
    43: T0 = 32'h3ffc28ac;
    44: T0 = 32'he8300002;
    45: T0 = 32'hffffe644;
    46: T0 = 32'hddbe2000;
    47: T0 = 32'h2f7a89ea;
    48: T0 = 32'h90a13ccb;
    49: T0 = 32'hd3f0f667;
    50: T0 = 32'hddaeecd6;
    51: T0 = 32'h71e35dec;
    52: T0 = 32'hfbdba171;
    53: T0 = 32'hee2b0142;
    54: T0 = 32'hb3800090;
    55: T0 = 32'hf95d000c;
    56: T0 = 32'h2007c06a;
    57: T0 = 32'h3fd288df;
    58: T0 = 32'ha700fe04;
    59: T0 = 32'hb7f2d45;
    60: T0 = 32'hfa407f80;
    61: T0 = 32'h807f03c0;
    62: T0 = 32'hc59145f0;
    63: T0 = 32'h201f0019;
    64: T0 = 32'he031f0ff;
    65: T0 = 32'h3c07f0c7;
    66: T0 = 32'h7e00fc87;
    67: T0 = 32'h7f03;
    68: T0 = 32'h7e07f90;
    69: T0 = 32'h374fe0;
    70: T0 = 32'hf07c071c;
    71: T0 = 32'hee08bddc;
    72: T0 = 32'h6b87c001;
    73: T0 = 32'h7ffcfafe;
    74: T0 = 32'h6987400;
    75: T0 = 32'h83f71f6f;
    76: T0 = 32'he18741c0;
    77: T0 = 32'hfc3907f5;
    78: T0 = 32'hc00afc2e;
    79: T0 = 32'h8f8061f2;
    80: T0 = 32'h4002000;
    81: T0 = 32'h5bc021e;
    82: T0 = 32'hd040cad4;
    83: T0 = 32'hd786f1;
    84: T0 = 32'ha3021c70;
    85: T0 = 32'h1edda7ff;
    86: T0 = 32'hd06ff0f4;
    87: T0 = 32'hff58bf;
    88: T0 = 32'hf740fe0f;
    89: T0 = 32'he07fadf;
    90: T0 = 32'h3f132ff0;
    91: T0 = 32'h4c2007f6;
    92: T0 = 32'h2d7002f8;
    93: T0 = 32'h39be907d;
    94: T0 = 32'h702f1d23;
    95: T0 = 32'h88d2c9e6;
    96: T0 = 32'h7e408f75;
    97: T0 = 32'h6a36849f;
    98: T0 = 32'hc885c7b8;
    99: T0 = 32'hbd8c1ddb;
    100: T0 = 32'h34855800;
    101: T0 = 32'h8b886e92;
    102: T0 = 32'hc7da8a76;
    103: T0 = 32'h1ccd7f9f;
    104: T0 = 32'hf5b60fe9;
    105: T0 = 32'h53c10acf;
    106: T0 = 32'h78209fe;
    107: T0 = 32'hd4ff83ef;
    108: T0 = 32'ha270049f;
    109: T0 = 32'h837ff870;
    110: T0 = 32'hf1e8c001;
    111: T0 = 32'hd00b2fc7;
    112: T0 = 32'h7f1f3e05;
    113: T0 = 32'h7d041ff8;
    114: T0 = 32'h37f0c1fc;
    115: T0 = 32'h81e4cd8f;
    116: T0 = 32'he1fffc1f;
    117: T0 = 32'hf81fff65;
    118: T0 = 32'h1c7377e0;
    119: T0 = 32'hafc001d9;
    120: T0 = 32'h3f8353f;
    121: T0 = 32'h75fef0cb;
    122: T0 = 32'hebcbff60;
    123: T0 = 32'h4149019e;
    124: T0 = 32'h13dd68e;
    125: T0 = 32'hfb52f010;
    126: T0 = 32'h60139e24;
    127: T0 = 32'h3e7cb103;
    128: T0 = 32'hcf82e1ed;
    129: T0 = 32'h83f5ff25;
    130: T0 = 32'hfff957df;
    131: T0 = 32'h803fff9d;
    132: T0 = 32'hf7d3dc01;
    133: T0 = 32'hac131f3f;
    134: T0 = 32'h1ffbc5c8;
    135: T0 = 32'hc9e007db;
    136: T0 = 32'h1ffe84f;
    137: T0 = 32'hff6e507b;
    138: T0 = 32'he01f5f07;
    139: T0 = 32'hfcf1b90f;
    140: T0 = 32'h8101b1fb;
    141: T0 = 32'h1c41ff89;
    142: T0 = 32'hb280fd6d;
    143: T0 = 32'hf4eafc23;
    144: T0 = 32'h31cd7ff3;
    145: T0 = 32'hcae06e2c;
    146: T0 = 32'h77beaa6b;
    147: T0 = 32'h5d27e3e0;
    148: T0 = 32'h4bb327ba;
    149: T0 = 32'hb64f13af;
    150: T0 = 32'hfc12ce57;
    151: T0 = 32'hf7f0fbb1;
    152: T0 = 32'h6c862e97;
    153: T0 = 32'h183c4b02;
    154: T0 = 32'hd4000d2b;
    155: T0 = 32'h2348718;
    156: T0 = 32'hdb60e7c0;
    157: T0 = 32'hc06c37df;
    158: T0 = 32'hfd9f0000;
    159: T0 = 32'hc4fd02e5;
    160: T0 = 32'hffcc6000;
    161: T0 = 32'h803f001a;
    162: T0 = 32'hff07c200;
    163: T0 = 32'ha010c05;
    164: T0 = 32'h5ffff890;
    165: T0 = 32'hbad883e1;
    166: T0 = 32'h7f7f9b;
    167: T0 = 32'h49e0f3f;
    168: T0 = 32'h5830fbe6;
    169: T0 = 32'h14704df;
    170: T0 = 32'h1de6ff17;
    171: T0 = 32'h44d5f;
    172: T0 = 32'hcdfcffe0;
    173: T0 = 32'he01701a3;
    174: T0 = 32'hd431ffc4;
    175: T0 = 32'h3f00401c;
    176: T0 = 32'h1d6088f8;
    177: T0 = 32'h2ff08601;
    178: T0 = 32'h81027afe;
    179: T0 = 32'h13386ff;
    180: T0 = 32'hfc00f4fc;
    181: T0 = 32'h35008f;
    182: T0 = 32'h26f0ffd5;
    183: T0 = 32'h1da07;
    184: T0 = 32'h890b3ffc;
    185: T0 = 32'hc0043f0;
    186: T0 = 32'he4d300c3;
    187: T0 = 32'h467a00bd;
    188: T0 = 32'hffdaf000;
    189: T0 = 32'h930f002c;
    190: T0 = 32'h7f88da40;
    191: T0 = 32'h83408000;
    192: T0 = 32'hfbf95e34;
    193: T0 = 32'h1db7402;
    194: T0 = 32'h7ffafd6d;
    195: T0 = 32'h76532fe6;
    196: T0 = 32'h64257b07;
    197: T0 = 32'h9cb41df2;
    198: T0 = 32'h10f8c4f1;
    199: T0 = 32'h5ffe3560;
    200: T0 = 32'ha37272a7;
    201: T0 = 32'hff046fdd;
    202: T0 = 32'ha3c9101c;
    203: T0 = 32'h13000151;
    204: T0 = 32'h19cb6200;
    205: T0 = 32'hc7a0c003;
    206: T0 = 32'h67dc2095;
    207: T0 = 32'hf9a03fc0;
    208: T0 = 32'hbfff0166;
    209: T0 = 32'hfd6e73ff;
    210: T0 = 32'hfffffc0d;
    211: T0 = 32'hff99abff;
    212: T0 = 32'hc3ff7fe1;
    213: T0 = 32'hf7fbad3f;
    214: T0 = 32'hfe7ffbff;
    215: T0 = 32'hfe3ff9c7;
    216: T0 = 32'hff24bffe;
    217: T0 = 32'hcfe3e09f;
    218: T0 = 32'h3ffd07d8;
    219: T0 = 32'h241e0403;
    220: T0 = 32'he3ff380c;
    221: T0 = 32'h27c12040;
    222: T0 = 32'he20032f;
    223: T0 = 32'hc8fc00;
    224: T0 = 32'hc0301105;
    225: T0 = 32'h3a800;
    226: T0 = 32'he7028002;
    227: T0 = 32'hf000c660;
    228: T0 = 32'h625f0e01;
    229: T0 = 32'h6d003690;
    230: T0 = 32'hff091e4;
    231: T0 = 32'hdf6423f8;
    232: T0 = 32'h60fad20c;
    233: T0 = 32'h9ff8081f;
    234: T0 = 32'h2bfd0c0;
    235: T0 = 32'hd3bf0142;
    236: T0 = 32'hf07fff68;
    237: T0 = 32'hf90ce202;
    238: T0 = 32'he2fffd8;
    239: T0 = 32'hfc08a066;
    240: T0 = 32'he03ffff2;
    241: T0 = 32'hffb3c02f;
    242: T0 = 32'hc1c2fffc;
    243: T0 = 32'h1b523970;
    244: T0 = 32'h981e3dd7;
    245: T0 = 32'hd5f43d26;
    246: T0 = 32'h133ee85b;
    247: T0 = 32'hedd138ea;
    248: T0 = 32'hff298018;
    249: T0 = 32'h97f1000a;
    250: T0 = 32'hfaf8030d;
    251: T0 = 32'hfc938000;
    252: T0 = 32'hd41f0013;
    253: T0 = 32'hffc70900;
    254: T0 = 32'h56890003;
    255: T0 = 32'h9fff11a8;
    256: T0 = 32'hef71b7f8;
    257: T0 = 32'h3fdf003;
    258: T0 = 32'hbbfeff;
    259: T0 = 32'ha0ffffd5;
    260: T0 = 32'hf003c7ef;
    261: T0 = 32'h2a1f7fec;
    262: T0 = 32'hfe407efe;
    263: T0 = 32'h183f7fe;
    264: T0 = 32'h3fc0dfdf;
    265: T0 = 32'h1038ffff;
    266: T0 = 32'hc3fc00bf;
    267: T0 = 32'hc3c7463e;
    268: T0 = 32'h4c1f2000;
    269: T0 = 32'hfe1c0940;
    270: T0 = 32'h61c01004;
    271: T0 = 32'h3e0c042;
    272: T0 = 32'h7a45940;
    273: T0 = 32'h1f0f0e;
    274: T0 = 32'h3619f57e;
    275: T0 = 32'h800039ff;
    276: T0 = 32'h3f3f073;
    277: T0 = 32'h3fc0008f;
    278: T0 = 32'hc0f1fa2;
    279: T0 = 32'h7fdc2be0;
    280: T0 = 32'hd84001f3;
    281: T0 = 32'hc4bddf98;
    282: T0 = 32'h8afc800f;
    283: T0 = 32'h23bfb6f0;
    284: T0 = 32'h7d7f4000;
    285: T0 = 32'hc075fd11;
    286: T0 = 32'h83e95800;
    287: T0 = 32'h507bffea;
    288: T0 = 32'hbdb95bc1;
    289: T0 = 32'h104fffff;
    290: T0 = 32'hff3c9087;
    291: T0 = 32'hbe07eff;
    292: T0 = 32'hc7f2dcf2;
    293: T0 = 32'hb352d110;
    294: T0 = 32'had360735;
    295: T0 = 32'h509aa46;
    296: T0 = 32'h85581a28;
    297: T0 = 32'h19ca62f8;
    298: T0 = 32'he17c7dd5;
    299: T0 = 32'he3d07cd5;
    300: T0 = 32'h2e0911d0;
    301: T0 = 32'h1200f07e;
    302: T0 = 32'h1d563b4f;
    303: T0 = 32'h2a60fcbf;
    304: T0 = 32'h636de7a1;
    305: T0 = 32'h79d53f07;
    306: T0 = 32'hf87f0310;
    307: T0 = 32'hbee3a7e0;
    308: T0 = 32'h7bfd000c;
    309: T0 = 32'hfeb773fe;
    310: T0 = 32'h69820000;
    311: T0 = 32'h40f1e7f;
    312: T0 = 32'h3400f03e;
    313: T0 = 32'hfa77;
    314: T0 = 32'h184ff03;
    315: T0 = 32'h3feb;
    316: T0 = 32'h78139bf0;
    317: T0 = 32'h560081fe;
    318: T0 = 32'h7e1ff7f;
    319: T0 = 32'hd280ff0f;
    320: T0 = 32'h773f67;
    321: T0 = 32'hfea4e7f1;
    322: T0 = 32'h710381ec;
    323: T0 = 32'h7c00469f;
    324: T0 = 32'h27e83c1f;
    325: T0 = 32'h4000f6cf;
    326: T0 = 32'h7dfc961;
    327: T0 = 32'hff001e63;
    328: T0 = 32'h121ece;
    329: T0 = 32'h8ff023f4;
    330: T0 = 32'h8005a6f4;
    331: T0 = 32'hadff533f;
    332: T0 = 32'hff0196ce;
    333: T0 = 32'hfeff3a5f;
    334: T0 = 32'hc47ff2ed;
    335: T0 = 32'hffd2f011;
    336: T0 = 32'h1c0feff2;
    337: T0 = 32'h7ff074bf;
    338: T0 = 32'hbbc288ff;
    339: T0 = 32'ha7ffe7ff;
    340: T0 = 32'h2efe181f;
    341: T0 = 32'h40193942;
    342: T0 = 32'h8a9b6bb0;
    343: T0 = 32'h71e7d6e7;
    344: T0 = 32'hed612cb1;
    345: T0 = 32'hb3796182;
    346: T0 = 32'hb9f7f997;
    347: T0 = 32'ha79d0c1e;
    348: T0 = 32'h8002794f;
    349: T0 = 32'h54d1500;
    350: T0 = 32'h2f6;
    351: T0 = 32'h902b1500;
    352: T0 = 32'h6900002f;
    353: T0 = 32'h283ad48;
    354: T0 = 32'he984001;
    355: T0 = 32'hce791e9b;
    356: T0 = 32'hd2ab6a00;
    357: T0 = 32'h3ff8037c;
    358: T0 = 32'hc6812a3e;
    359: T0 = 32'h1bfffca0;
    360: T0 = 32'hf8ea03f7;
    361: T0 = 32'hec3f7fd0;
    362: T0 = 32'hef1fea77;
    363: T0 = 32'hfedfbe78;
    364: T0 = 32'h3f018464;
    365: T0 = 32'h3ff2c9d5;
    366: T0 = 32'ha078e841;
    367: T0 = 32'hc3fff31f;
    368: T0 = 32'hfbc7ff85;
    369: T0 = 32'he1f1bab;
    370: T0 = 32'hff2a1ffc;
    371: T0 = 32'h61e3fc;
    372: T0 = 32'h7f3076f;
    373: T0 = 32'h70037f3f;
    374: T0 = 32'h32776bc9;
    375: T0 = 32'he5a003fe;
    376: T0 = 32'ha21f2f2;
    377: T0 = 32'h1e58a007;
    378: T0 = 32'h45830002;
    379: T0 = 32'h10c3a600;
    380: T0 = 32'h4c330000;
    381: T0 = 32'h118206b0;
    382: T0 = 32'h39f0000;
    383: T0 = 32'hf72203cf;
    384: T0 = 32'h174000;
    385: T0 = 32'h17fc003c;
    386: T0 = 32'h8008d200;
    387: T0 = 32'hfbfbf028;
    388: T0 = 32'hc0049a4e;
    389: T0 = 32'h3685a580;
    390: T0 = 32'h376db407;
    391: T0 = 32'hedefc7a0;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T5 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T6 = reset ? 1'h0 : restartRegs_0;
  assign T7 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_3(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T5;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T6;
  reg  restartRegs_0;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (addr)
    0: T0 = 32'ha3cfbde;
    1: T0 = 32'h7759acd2;
    2: T0 = 32'h40e26470;
    3: T0 = 32'h700759fe;
    4: T0 = 32'h16cba4b8;
    5: T0 = 32'h227ab687;
    6: T0 = 32'hf96de001;
    7: T0 = 32'h68170009;
    8: T0 = 32'hbfee0b80;
    9: T0 = 32'h4cf0a70c;
    10: T0 = 32'h1ff63299;
    11: T0 = 32'he0673ac0;
    12: T0 = 32'hb81f0697;
    13: T0 = 32'hfe24ff90;
    14: T0 = 32'ha3800037;
    15: T0 = 32'hff7efbd;
    16: T0 = 32'h3a1c8080;
    17: T0 = 32'he17e0b3d;
    18: T0 = 32'hf947f80e;
    19: T0 = 32'hff03f057;
    20: T0 = 32'hf617ecf;
    21: T0 = 32'h1ff8ff01;
    22: T0 = 32'h80fa2b81;
    23: T0 = 32'h85ff3ff0;
    24: T0 = 32'hd2070090;
    25: T0 = 32'hf87f01ff;
    26: T0 = 32'hf9b0e059;
    27: T0 = 32'hf5b383f;
    28: T0 = 32'hff8ff803;
    29: T0 = 32'hb0c41f03;
    30: T0 = 32'h7f783b00;
    31: T0 = 32'hd3bc6090;
    32: T0 = 32'h8bff03e0;
    33: T0 = 32'hff1f1233;
    34: T0 = 32'hf9c0f03e;
    35: T0 = 32'he7e0cf48;
    36: T0 = 32'h87fd9f83;
    37: T0 = 32'h467c39cf;
    38: T0 = 32'h803ffb58;
    39: T0 = 32'hfb8f00bf;
    40: T0 = 32'hfdfbb26b;
    41: T0 = 32'h1fba101f;
    42: T0 = 32'h79ea803;
    43: T0 = 32'h36fea083;
    44: T0 = 32'hb2f94000;
    45: T0 = 32'h8a8f1340;
    46: T0 = 32'h7873d20;
    47: T0 = 32'h3008385a;
    48: T0 = 32'h643cd8ed;
    49: T0 = 32'h8d52ab9a;
    50: T0 = 32'h541f9abf;
    51: T0 = 32'h8a20c299;
    52: T0 = 32'h72e708b8;
    53: T0 = 32'hca6fffbb;
    54: T0 = 32'h74407c00;
    55: T0 = 32'he91e7ffe;
    56: T0 = 32'h636c64ac;
    57: T0 = 32'h7fe8c9fe;
    58: T0 = 32'h8e3ce132;
    59: T0 = 32'h8fff369f;
    60: T0 = 32'hf718dff4;
    61: T0 = 32'h57ff002e;
    62: T0 = 32'hafe4b01c;
    63: T0 = 32'ha1bf0002;
    64: T0 = 32'hf8f15840;
    65: T0 = 32'h8c5f0000;
    66: T0 = 32'hfe0780c0;
    67: T0 = 32'h17031000;
    68: T0 = 32'hffc05760;
    69: T0 = 32'h30447d0;
    70: T0 = 32'h1ff8fff9;
    71: T0 = 32'h1e81ef;
    72: T0 = 32'hb1ffffff;
    73: T0 = 32'he003fe7e;
    74: T0 = 32'hf89e4fff;
    75: T0 = 32'hfe0affb7;
    76: T0 = 32'h7e6d8bbf;
    77: T0 = 32'h1ff0fbf8;
    78: T0 = 32'h3e1b80f;
    79: T0 = 32'hf5fffe0d;
    80: T0 = 32'hf80f1185;
    81: T0 = 32'hf4d77fc0;
    82: T0 = 32'h3f8001fa;
    83: T0 = 32'h3ca07f0;
    84: T0 = 32'h40e40019;
    85: T0 = 32'h3f667e;
    86: T0 = 32'hd400e680;
    87: T0 = 32'hd83040f;
    88: T0 = 32'h83407c00;
    89: T0 = 32'h81910fd6;
    90: T0 = 32'hfa1f4fc0;
    91: T0 = 32'h1c223fec;
    92: T0 = 32'hd0da79ed;
    93: T0 = 32'h1ac23fff;
    94: T0 = 32'hbfff563;
    95: T0 = 32'h92a02677;
    96: T0 = 32'h973b509b;
    97: T0 = 32'hdf020ec0;
    98: T0 = 32'h2dae0292;
    99: T0 = 32'hab13890e;
    100: T0 = 32'h6ffdb3fb;
    101: T0 = 32'hbb8ec756;
    102: T0 = 32'hcf80c5f2;
    103: T0 = 32'h6db5b052;
    104: T0 = 32'h2866f826;
    105: T0 = 32'h3fe06238;
    106: T0 = 32'h80382aba;
    107: T0 = 32'h2fff6f09;
    108: T0 = 32'hff680628;
    109: T0 = 32'ha77900c3;
    110: T0 = 32'h800d1454;
    111: T0 = 32'h3e987807;
    112: T0 = 32'hf800f2a3;
    113: T0 = 32'h5ef43fb;
    114: T0 = 32'h4400e705;
    115: T0 = 32'h7fc87f;
    116: T0 = 32'hf582fc24;
    117: T0 = 32'h207064f;
    118: T0 = 32'hff58ff80;
    119: T0 = 32'he10074;
    120: T0 = 32'h1faa67f8;
    121: T0 = 32'hbde60065;
    122: T0 = 32'he1e4c6ff;
    123: T0 = 32'he59c904f;
    124: T0 = 32'he71efc1a;
    125: T0 = 32'h9e07810f;
    126: T0 = 32'h2d2f7fe4;
    127: T0 = 32'hf82f4e00;
    128: T0 = 32'h68010ff2;
    129: T0 = 32'h87c084b6;
    130: T0 = 32'ha20307f;
    131: T0 = 32'h33ee84b;
    132: T0 = 32'he0d5cf07;
    133: T0 = 32'hfb7ffe83;
    134: T0 = 32'hfe0a0ee0;
    135: T0 = 32'heb4607ed;
    136: T0 = 32'h7fe0f7de;
    137: T0 = 32'h22ce07f;
    138: T0 = 32'h3fbcff8f;
    139: T0 = 32'h30e9e01;
    140: T0 = 32'ha7ee1fe1;
    141: T0 = 32'h325660;
    142: T0 = 32'h9e28005c;
    143: T0 = 32'hfab98;
    144: T0 = 32'hf420a525;
    145: T0 = 32'h41000721;
    146: T0 = 32'heb9ee7db;
    147: T0 = 32'h97a6c4ea;
    148: T0 = 32'h461c910a;
    149: T0 = 32'hd02661aa;
    150: T0 = 32'h1e19ce96;
    151: T0 = 32'h5f124bf0;
    152: T0 = 32'h1e0115b;
    153: T0 = 32'h88c0a617;
    154: T0 = 32'h803f04a9;
    155: T0 = 32'h7db670b7;
    156: T0 = 32'h66000125;
    157: T0 = 32'h1ff32ffe;
    158: T0 = 32'h681ce84d;
    159: T0 = 32'hc07ef053;
    160: T0 = 32'hc5c77ff5;
    161: T0 = 32'h3e03fdff;
    162: T0 = 32'h3d482bff;
    163: T0 = 32'h1ff0fe98;
    164: T0 = 32'h23e30bdb;
    165: T0 = 32'h3e7f01e0;
    166: T0 = 32'h423c2c29;
    167: T0 = 32'he70000;
    168: T0 = 32'h70310153;
    169: T0 = 32'h72090800;
    170: T0 = 32'h2e060001;
    171: T0 = 32'h7fe00a80;
    172: T0 = 32'h0;
    173: T0 = 32'h7380028;
    174: T0 = 32'hc054c006;
    175: T0 = 32'h607f7001;
    176: T0 = 32'h7c015800;
    177: T0 = 32'hcb070fc0;
    178: T0 = 32'h738519c0;
    179: T0 = 32'h7f3203fc;
    180: T0 = 32'hc39dba0c;
    181: T0 = 32'h79c7687f;
    182: T0 = 32'h9e78ffde;
    183: T0 = 32'h83cbdbbf;
    184: T0 = 32'h68effe1e;
    185: T0 = 32'hf83fbb4c;
    186: T0 = 32'hf3bf9fc4;
    187: T0 = 32'h8f81fe55;
    188: T0 = 32'h9fd0efbb;
    189: T0 = 32'h90f8dfa8;
    190: T0 = 32'h80fc3cbe;
    191: T0 = 32'h9f0fcffb;
    192: T0 = 32'hf8074aab;
    193: T0 = 32'h2a903fdd;
    194: T0 = 32'h8f80a5a3;
    195: T0 = 32'h50c13db7;
    196: T0 = 32'hd15e87a;
    197: T0 = 32'hb977e0e;
    198: T0 = 32'hdb99f0b1;
    199: T0 = 32'h9133f840;
    200: T0 = 32'h95c2efd8;
    201: T0 = 32'h18112b8;
    202: T0 = 32'h1c87860;
    203: T0 = 32'h57300001;
    204: T0 = 32'h5eec47;
    205: T0 = 32'h7738f001;
    206: T0 = 32'haa0211f1;
    207: T0 = 32'h15d07c00;
    208: T0 = 32'h1f60045e;
    209: T0 = 32'h5fe6c0;
    210: T0 = 32'hf9a81bfe;
    211: T0 = 32'hc023b038;
    212: T0 = 32'h2721fffe;
    213: T0 = 32'h7e02fe3f;
    214: T0 = 32'h66fefdff;
    215: T0 = 32'hc9e0ffe7;
    216: T0 = 32'h8bdfb307;
    217: T0 = 32'hf01f3fbd;
    218: T0 = 32'hfc3eee40;
    219: T0 = 32'h4e000017;
    220: T0 = 32'h7c10df8;
    221: T0 = 32'h3040c000;
    222: T0 = 32'h41e20f9;
    223: T0 = 32'h3c85200;
    224: T0 = 32'hc1c18298;
    225: T0 = 32'h282fef;
    226: T0 = 32'hac0e7811;
    227: T0 = 32'he007b13c;
    228: T0 = 32'hfb80efc1;
    229: T0 = 32'hfe03f73;
    230: T0 = 32'hffca1ed2;
    231: T0 = 32'h607f03d2;
    232: T0 = 32'hfd5f8800;
    233: T0 = 32'hf803007d;
    234: T0 = 32'h3ff155a0;
    235: T0 = 32'hde08007;
    236: T0 = 32'h1e2ffcf;
    237: T0 = 32'hf9ba1049;
    238: T0 = 32'h74014a5b;
    239: T0 = 32'h75159f;
    240: T0 = 32'h41f0ff83;
    241: T0 = 32'h40175e98;
    242: T0 = 32'h91f9093;
    243: T0 = 32'h27110d70;
    244: T0 = 32'hc22ae9d1;
    245: T0 = 32'h9bbfff0a;
    246: T0 = 32'h544a0ca1;
    247: T0 = 32'h4bc0e47e;
    248: T0 = 32'ha0366c75;
    249: T0 = 32'h68a9b78b;
    250: T0 = 32'hfffefa56;
    251: T0 = 32'hcb84e834;
    252: T0 = 32'h19ff0acc;
    253: T0 = 32'h3a525436;
    254: T0 = 32'hd20ef178;
    255: T0 = 32'h174016f;
    256: T0 = 32'h8240f81e;
    257: T0 = 32'h3d1f86d;
    258: T0 = 32'hdef13e40;
    259: T0 = 32'hd03f1fc6;
    260: T0 = 32'he1fe2be0;
    261: T0 = 32'hd7c101f8;
    262: T0 = 32'hf9389fc;
    263: T0 = 32'hfc6ec01f;
    264: T0 = 32'hf077f879;
    265: T0 = 32'h7f2c5801;
    266: T0 = 32'h6fc03c00;
    267: T0 = 32'h1b845c4;
    268: T0 = 32'h63fe03e0;
    269: T0 = 32'hf82384bf;
    270: T0 = 32'h1fff503f;
    271: T0 = 32'hffc0fcd9;
    272: T0 = 32'h48ad203;
    273: T0 = 32'h57fc3ffd;
    274: T0 = 32'hf0003b8c;
    275: T0 = 32'h9813c3ff;
    276: T0 = 32'h9f80f4b3;
    277: T0 = 32'h7c0c51f;
    278: T0 = 32'hf8fb7b;
    279: T0 = 32'h85681e09;
    280: T0 = 32'hc02f1f80;
    281: T0 = 32'hf80c6380;
    282: T0 = 32'hd80201ff;
    283: T0 = 32'h6f84c33f;
    284: T0 = 32'h820001d;
    285: T0 = 32'hc01f0b7;
    286: T0 = 32'h53a01b;
    287: T0 = 32'habf0b814;
    288: T0 = 32'hc0dee801;
    289: T0 = 32'he1f90000;
    290: T0 = 32'hdd9f2a34;
    291: T0 = 32'h35f4e04;
    292: T0 = 32'hc7ffa226;
    293: T0 = 32'h2ca367bc;
    294: T0 = 32'h24fb399c;
    295: T0 = 32'h80b2ed21;
    296: T0 = 32'h92aecd6e;
    297: T0 = 32'h742805c8;
    298: T0 = 32'h39549832;
    299: T0 = 32'h6bc42f75;
    300: T0 = 32'h1300b7f;
    301: T0 = 32'he200cd8e;
    302: T0 = 32'hde8648;
    303: T0 = 32'h52e02429;
    304: T0 = 32'h4038068;
    305: T0 = 32'hcd81d7f;
    306: T0 = 32'h1ffcfc9a;
    307: T0 = 32'hfde8807f;
    308: T0 = 32'h87ffff46;
    309: T0 = 32'hffd940a3;
    310: T0 = 32'h6caf8140;
    311: T0 = 32'hfffe07c0;
    312: T0 = 32'hea9cc000;
    313: T0 = 32'hc0ff801d;
    314: T0 = 32'h7faffe73;
    315: T0 = 32'h5fcefc00;
    316: T0 = 32'hc01957ff;
    317: T0 = 32'h7ffefffc;
    318: T0 = 32'h9c01e07f;
    319: T0 = 32'hee3ffbf;
    320: T0 = 32'h40e0ff77;
    321: T0 = 32'h3a3ff9;
    322: T0 = 32'hd0060ffb;
    323: T0 = 32'h350083ff;
    324: T0 = 32'h6c00e0ff;
    325: T0 = 32'h774fd3f;
    326: T0 = 32'ha5b0f807;
    327: T0 = 32'h906f1f27;
    328: T0 = 32'h41f7e00;
    329: T0 = 32'hfe800022;
    330: T0 = 32'hc1fea0;
    331: T0 = 32'h39f80000;
    332: T0 = 32'hf0144f2c;
    333: T0 = 32'h66bf0024;
    334: T0 = 32'h9fef1d66;
    335: T0 = 32'hfdc6f000;
    336: T0 = 32'h8ff0cf0;
    337: T0 = 32'hffeba090;
    338: T0 = 32'hdae73f9d;
    339: T0 = 32'hfffa4243;
    340: T0 = 32'h67fb34e0;
    341: T0 = 32'h3fffe914;
    342: T0 = 32'h66e3cc82;
    343: T0 = 32'ha9ed8cac;
    344: T0 = 32'hfd7596ab;
    345: T0 = 32'h6211f1ca;
    346: T0 = 32'hae5c4f2e;
    347: T0 = 32'heb5699ed;
    348: T0 = 32'h7fdaed2f;
    349: T0 = 32'hfea6e98f;
    350: T0 = 32'he3ffffda;
    351: T0 = 32'he663f31f;
    352: T0 = 32'he50f5ff9;
    353: T0 = 32'h304f0;
    354: T0 = 32'hd2000ffc;
    355: T0 = 32'ha002e;
    356: T0 = 32'hfa4ce1fe;
    357: T0 = 32'hc000c004;
    358: T0 = 32'hfdfee43f;
    359: T0 = 32'hc00f800;
    360: T0 = 32'h1fff06a7;
    361: T0 = 32'h3fc87f00;
    362: T0 = 32'h80f5038e;
    363: T0 = 32'h2bd8c7e0;
    364: T0 = 32'h1f5f023b;
    365: T0 = 32'h1fbd07e;
    366: T0 = 32'hf5e7a053;
    367: T0 = 32'h7001bfa3;
    368: T0 = 32'h7e1f01;
    369: T0 = 32'hfe005fd8;
    370: T0 = 32'h638060;
    371: T0 = 32'h3fcc0531;
    372: T0 = 32'he087f002;
    373: T0 = 32'h6ffc1013;
    374: T0 = 32'h5e083d40;
    375: T0 = 32'hcb309d6;
    376: T0 = 32'hc6f89762;
    377: T0 = 32'h8005f1ff;
    378: T0 = 32'hcedf3e72;
    379: T0 = 32'hfc3cd1ef;
    380: T0 = 32'hf60fd02b;
    381: T0 = 32'h7fc08e8e;
    382: T0 = 32'h15801f9f;
    383: T0 = 32'h184fcf;
    384: T0 = 32'h40bdf3ea;
    385: T0 = 32'hf000b7ec;
    386: T0 = 32'h7519c4f9;
    387: T0 = 32'hd80e1f8;
    388: T0 = 32'hff9feffd;
    389: T0 = 32'h9e60ae0f;
    390: T0 = 32'h4f363c00;
    391: T0 = 32'h8fa6d1fc;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T5 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T6 = reset ? 1'h0 : restartRegs_0;
  assign T7 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_4(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T5;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T6;
  reg  restartRegs_0;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (addr)
    0: T0 = 32'h9a165153;
    1: T0 = 32'h83e25630;
    2: T0 = 32'hd475459b;
    3: T0 = 32'h6705c0f8;
    4: T0 = 32'hf6c5bf91;
    5: T0 = 32'hf44c0a8d;
    6: T0 = 32'h9cdec5fe;
    7: T0 = 32'h88800fd;
    8: T0 = 32'had29de;
    9: T0 = 32'h27f1c00c;
    10: T0 = 32'h1002ad87;
    11: T0 = 32'hc5bc0003;
    12: T0 = 32'hf8007c0;
    13: T0 = 32'h1dd000c0;
    14: T0 = 32'hc1fc0376;
    15: T0 = 32'hc3f7c007;
    16: T0 = 32'hcc0f1c0f;
    17: T0 = 32'h7c3d16c0;
    18: T0 = 32'hda400970;
    19: T0 = 32'h7c7c3b8;
    20: T0 = 32'h7ea681f3;
    21: T0 = 32'hc17c9e0a;
    22: T0 = 32'hc7f8603d;
    23: T0 = 32'h9297e9f0;
    24: T0 = 32'hfc2e1903;
    25: T0 = 32'hffd73f0f;
    26: T0 = 32'hffc2f0e4;
    27: T0 = 32'h37c703f9;
    28: T0 = 32'h63f89f04;
    29: T0 = 32'h8fff81f;
    30: T0 = 32'h984ffcf0;
    31: T0 = 32'h1b500b03;
    32: T0 = 32'h2007ce;
    33: T0 = 32'h308028;
    34: T0 = 32'h78c3af;
    35: T0 = 32'hc000f013;
    36: T0 = 32'h70290;
    37: T0 = 32'hcc00ef03;
    38: T0 = 32'h753c;
    39: T0 = 32'h78ccc3f0;
    40: T0 = 32'hc00cc162;
    41: T0 = 32'h7fe5c9c9;
    42: T0 = 32'hb000bc0c;
    43: T0 = 32'ha7fb8df7;
    44: T0 = 32'h663e1fc0;
    45: T0 = 32'hffff3015;
    46: T0 = 32'hf7c147fe;
    47: T0 = 32'ha13f1d0f;
    48: T0 = 32'h207071f;
    49: T0 = 32'hc6c66546;
    50: T0 = 32'h5e953034;
    51: T0 = 32'h350c666b;
    52: T0 = 32'hbb92ed2b;
    53: T0 = 32'h2d153bb1;
    54: T0 = 32'hd9743057;
    55: T0 = 32'he34bc43b;
    56: T0 = 32'h137f806e;
    57: T0 = 32'h5d2bac17;
    58: T0 = 32'h30ff001;
    59: T0 = 32'hfff10fa0;
    60: T0 = 32'h5b37f03;
    61: T0 = 32'hf9c27f94;
    62: T0 = 32'h9303e0;
    63: T0 = 32'h3efc0ffe;
    64: T0 = 32'h1644ae3f;
    65: T0 = 32'h9079f8ff;
    66: T0 = 32'h1e0f9a0;
    67: T0 = 32'h17000f83;
    68: T0 = 32'h21f0621;
    69: T0 = 32'hc1488078;
    70: T0 = 32'h80ffc038;
    71: T0 = 32'hfc080687;
    72: T0 = 32'hea07b801;
    73: T0 = 32'hff8000df;
    74: T0 = 32'h6f0ffd0;
    75: T0 = 32'h2f0c079;
    76: T0 = 32'h1d75fdd;
    77: T0 = 32'he507e33f;
    78: T0 = 32'h8012ed3f;
    79: T0 = 32'hfc31e683;
    80: T0 = 32'hf8073940;
    81: T0 = 32'h7fe30210;
    82: T0 = 32'h3b800b92;
    83: T0 = 32'hfeaa002;
    84: T0 = 32'h21988dbb;
    85: T0 = 32'hc7f1b500;
    86: T0 = 32'h3d0b0f7c;
    87: T0 = 32'h22fbf1c0;
    88: T0 = 32'h801001c3;
    89: T0 = 32'h1fc0ffe;
    90: T0 = 32'hffdf701b;
    91: T0 = 32'h701f9afd;
    92: T0 = 32'h7ff21383;
    93: T0 = 32'heb002710;
    94: T0 = 32'hfea230;
    95: T0 = 32'hd192bd01;
    96: T0 = 32'h8a9fe26f;
    97: T0 = 32'h8b9bf7f3;
    98: T0 = 32'h60581d32;
    99: T0 = 32'h2fd544bb;
    100: T0 = 32'ha5356a1c;
    101: T0 = 32'h4f37239a;
    102: T0 = 32'h7bcec602;
    103: T0 = 32'h7f0000a5;
    104: T0 = 32'h3710140;
    105: T0 = 32'h9fe0e03e;
    106: T0 = 32'h71fe0f;
    107: T0 = 32'hc5fcff00;
    108: T0 = 32'h40313333;
    109: T0 = 32'h1cbf3f80;
    110: T0 = 32'hf000f6b2;
    111: T0 = 32'h1f743e1;
    112: T0 = 32'h3d001bed;
    113: T0 = 32'hff47e;
    114: T0 = 32'hab00e077;
    115: T0 = 32'h2bf1e07;
    116: T0 = 32'hfc80ff00;
    117: T0 = 32'hff6fc8;
    118: T0 = 32'hffd40ff0;
    119: T0 = 32'h807f00b8;
    120: T0 = 32'hfffaa3ff;
    121: T0 = 32'hfc17f877;
    122: T0 = 32'h7efff3bf;
    123: T0 = 32'h3651ffc0;
    124: T0 = 32'hcf433f64;
    125: T0 = 32'hb09787fe;
    126: T0 = 32'hd5e5f3f0;
    127: T0 = 32'h7804e04b;
    128: T0 = 32'he9fe1ffb;
    129: T0 = 32'hc600bb40;
    130: T0 = 32'hedf00f7;
    131: T0 = 32'hfcf13d82;
    132: T0 = 32'h1af4008;
    133: T0 = 32'h8fef00e7;
    134: T0 = 32'h68179000;
    135: T0 = 32'he2ff0f7f;
    136: T0 = 32'hde70e710;
    137: T0 = 32'h31eb00ff;
    138: T0 = 32'hff400815;
    139: T0 = 32'h63f881e;
    140: T0 = 32'h3ff0febb;
    141: T0 = 32'h8642c43;
    142: T0 = 32'h89dd1e21;
    143: T0 = 32'he002f020;
    144: T0 = 32'h383fef91;
    145: T0 = 32'hff845088;
    146: T0 = 32'hda507453;
    147: T0 = 32'hbfd9ff5d;
    148: T0 = 32'hfa510bc0;
    149: T0 = 32'h62cff065;
    150: T0 = 32'he288008e;
    151: T0 = 32'hacdf177;
    152: T0 = 32'h68cef9b;
    153: T0 = 32'hfea1419f;
    154: T0 = 32'he7ffffe1;
    155: T0 = 32'hd9caa71f;
    156: T0 = 32'hedf9cffc;
    157: T0 = 32'hdcb1fd43;
    158: T0 = 32'h99f01ff;
    159: T0 = 32'h24528222;
    160: T0 = 32'h80ae781f;
    161: T0 = 32'h100f804;
    162: T0 = 32'h7d132ffd;
    163: T0 = 32'h7c38fe00;
    164: T0 = 32'hff0f00ff;
    165: T0 = 32'h9d81ffc0;
    166: T0 = 32'h2ff200cf;
    167: T0 = 32'h4ece1fc;
    168: T0 = 32'hbffe005;
    169: T0 = 32'h3eec0b;
    170: T0 = 32'hf203df00;
    171: T0 = 32'h38a80;
    172: T0 = 32'h18f807f3;
    173: T0 = 32'hf40097fc;
    174: T0 = 32'h79f401f;
    175: T0 = 32'hfe0707a;
    176: T0 = 32'h1fbaf00;
    177: T0 = 32'hea7ca007;
    178: T0 = 32'h907fe073;
    179: T0 = 32'hfcafecc1;
    180: T0 = 32'hbfff1931;
    181: T0 = 32'hffc61ff8;
    182: T0 = 32'hf80f03f0;
    183: T0 = 32'h7ff20bfc;
    184: T0 = 32'h6db12043;
    185: T0 = 32'hb7e05bff;
    186: T0 = 32'h214a105;
    187: T0 = 32'hf34a087c;
    188: T0 = 32'h202afc00;
    189: T0 = 32'hb20894fa;
    190: T0 = 32'hd3e8ad42;
    191: T0 = 32'h9984ffea;
    192: T0 = 32'h4823e90b;
    193: T0 = 32'h64537ffa;
    194: T0 = 32'h20be1d8f;
    195: T0 = 32'h3a8159bb;
    196: T0 = 32'h3d872511;
    197: T0 = 32'hf71aba61;
    198: T0 = 32'hb1d749b5;
    199: T0 = 32'hc17f62de;
    200: T0 = 32'hef9ed7fd;
    201: T0 = 32'ha41afed7;
    202: T0 = 32'hf3f472ff;
    203: T0 = 32'he4c1f08b;
    204: T0 = 32'hf2af43f;
    205: T0 = 32'h5bf7fb08;
    206: T0 = 32'hf0e91421;
    207: T0 = 32'hced44000;
    208: T0 = 32'h2f0101f0;
    209: T0 = 32'h7ec49c00;
    210: T0 = 32'hc3e00000;
    211: T0 = 32'hfecf5fa;
    212: T0 = 32'h7aefe004;
    213: T0 = 32'hf87b5fff;
    214: T0 = 32'h783fffff;
    215: T0 = 32'hffc3ffef;
    216: T0 = 32'h5ff7fdf;
    217: T0 = 32'h5ffefffb;
    218: T0 = 32'hf0126829;
    219: T0 = 32'h2b31bfff;
    220: T0 = 32'hf80ba4a;
    221: T0 = 32'hef20bf8;
    222: T0 = 32'h23fe3fa8;
    223: T0 = 32'h8045807e;
    224: T0 = 32'h700fffb2;
    225: T0 = 32'hfa9c5803;
    226: T0 = 32'hfbbd1ffe;
    227: T0 = 32'h1fbfeb00;
    228: T0 = 32'hdd14c0ff;
    229: T0 = 32'hd67efef7;
    230: T0 = 32'he78fedb7;
    231: T0 = 32'he7431fd7;
    232: T0 = 32'h3d9041fe;
    233: T0 = 32'hed94e03c;
    234: T0 = 32'h41ef4f1e;
    235: T0 = 32'h57f8cc00;
    236: T0 = 32'h400f0b1b;
    237: T0 = 32'hfddc89e0;
    238: T0 = 32'ha0d8d06d;
    239: T0 = 32'h3f9e64b;
    240: T0 = 32'hf301f00f;
    241: T0 = 32'h87fe537;
    242: T0 = 32'hf8005beb;
    243: T0 = 32'h20217081;
    244: T0 = 32'h46111de;
    245: T0 = 32'h83a1ebf3;
    246: T0 = 32'ha5963f96;
    247: T0 = 32'h8aba0b87;
    248: T0 = 32'hde7c972d;
    249: T0 = 32'h9cdbfe1;
    250: T0 = 32'h5fe248c2;
    251: T0 = 32'he19cd23c;
    252: T0 = 32'h9effbf0f;
    253: T0 = 32'h7fd5c447;
    254: T0 = 32'h41fdf160;
    255: T0 = 32'hd41860ff;
    256: T0 = 32'h41d5ffc7;
    257: T0 = 32'hf4b08ad1;
    258: T0 = 32'hb383f9;
    259: T0 = 32'hf19c7961;
    260: T0 = 32'h12000;
    261: T0 = 32'hbf0000d7;
    262: T0 = 32'hb200;
    263: T0 = 32'h458000f1;
    264: T0 = 32'h900080a8;
    265: T0 = 32'h3bbc007f;
    266: T0 = 32'h9f80ff22;
    267: T0 = 32'hfff9140f;
    268: T0 = 32'hdeffff89;
    269: T0 = 32'hdfff13c1;
    270: T0 = 32'hf8477fe0;
    271: T0 = 32'h1ff014d;
    272: T0 = 32'hff085ff8;
    273: T0 = 32'h401f0011;
    274: T0 = 32'hffe0cdfe;
    275: T0 = 32'h4641c003;
    276: T0 = 32'hffc7def;
    277: T0 = 32'h8dc0f800;
    278: T0 = 32'h6ffc0fe0;
    279: T0 = 32'h232bf0e;
    280: T0 = 32'h4bf85ffa;
    281: T0 = 32'h804b2cd2;
    282: T0 = 32'hf3ff07ff;
    283: T0 = 32'hb2003c4b;
    284: T0 = 32'h33f0934;
    285: T0 = 32'hfe00e17a;
    286: T0 = 32'h73d83f9b;
    287: T0 = 32'h2ff062ea;
    288: T0 = 32'hfff28dc5;
    289: T0 = 32'h22ff1e0f;
    290: T0 = 32'hd778380d;
    291: T0 = 32'hed97e57f;
    292: T0 = 32'h275e7531;
    293: T0 = 32'ha0eb2043;
    294: T0 = 32'h4fab6c33;
    295: T0 = 32'h6bb8e8e8;
    296: T0 = 32'hf9b65091;
    297: T0 = 32'hf35a5bde;
    298: T0 = 32'he04ca6b1;
    299: T0 = 32'hbfc2c36a;
    300: T0 = 32'hd6dc35fd;
    301: T0 = 32'h2fe8ffdc;
    302: T0 = 32'h5fce6bb;
    303: T0 = 32'hdff9f9ff;
    304: T0 = 32'hcc1fb283;
    305: T0 = 32'h5ff0fff;
    306: T0 = 32'hc03f3ef4;
    307: T0 = 32'hf95d036e;
    308: T0 = 32'h5e0087f8;
    309: T0 = 32'h3b98020;
    310: T0 = 32'h3b007c3f;
    311: T0 = 32'h1ddfe80;
    312: T0 = 32'heb002fc3;
    313: T0 = 32'h3d3fd0;
    314: T0 = 32'hffb84160;
    315: T0 = 32'h783f03fe;
    316: T0 = 32'hbff39e9c;
    317: T0 = 32'he3ffe03f;
    318: T0 = 32'hf1fef7fe;
    319: T0 = 32'h44fffc0f;
    320: T0 = 32'hff1ffdfc;
    321: T0 = 32'he8438fc0;
    322: T0 = 32'h4ff11f81;
    323: T0 = 32'hef847ffe;
    324: T0 = 32'h383ee3f8;
    325: T0 = 32'hc780395f;
    326: T0 = 32'h783ff1e;
    327: T0 = 32'h3c39e7e8;
    328: T0 = 32'h12a01ff1;
    329: T0 = 32'h81e3b1f8;
    330: T0 = 32'h302ccc7f;
    331: T0 = 32'hd83efc03;
    332: T0 = 32'hf3d13567;
    333: T0 = 32'h3b017fc0;
    334: T0 = 32'hc7c03459;
    335: T0 = 32'h86d60ff8;
    336: T0 = 32'h7fee005;
    337: T0 = 32'hfc15c77f;
    338: T0 = 32'h827df807;
    339: T0 = 32'hc4138b8f;
    340: T0 = 32'hd857effa;
    341: T0 = 32'hbc0a737a;
    342: T0 = 32'h2c60e67c;
    343: T0 = 32'hb04f7081;
    344: T0 = 32'h496d775c;
    345: T0 = 32'h67a8d1a6;
    346: T0 = 32'hf977095f;
    347: T0 = 32'h24aa6c06;
    348: T0 = 32'he11877b0;
    349: T0 = 32'h7942bfe0;
    350: T0 = 32'hed105ffd;
    351: T0 = 32'hde5af2db;
    352: T0 = 32'h946f202f;
    353: T0 = 32'hf82248fc;
    354: T0 = 32'h25878080;
    355: T0 = 32'h3fe7009a;
    356: T0 = 32'h6a7fe000;
    357: T0 = 32'h35e50000;
    358: T0 = 32'h558c1800;
    359: T0 = 32'h43ef0140;
    360: T0 = 32'hfcc57700;
    361: T0 = 32'h25ff0006;
    362: T0 = 32'hf1f01ff8;
    363: T0 = 32'h1bf8040;
    364: T0 = 32'h7c0f03f8;
    365: T0 = 32'hf00d5a3c;
    366: T0 = 32'h3380f9ff;
    367: T0 = 32'h7f4d5e5;
    368: T0 = 32'h350afff;
    369: T0 = 32'h803ffd85;
    370: T0 = 32'hf61732ff;
    371: T0 = 32'h7a01ff8f;
    372: T0 = 32'hf9fe1ef;
    373: T0 = 32'h5ff87ff8;
    374: T0 = 32'ha07e61ff;
    375: T0 = 32'hf57fffff;
    376: T0 = 32'hff0783af;
    377: T0 = 32'h7f937ffc;
    378: T0 = 32'hdff0c0c8;
    379: T0 = 32'h87fa3dff;
    380: T0 = 32'he8fc031b;
    381: T0 = 32'he0ff32ee;
    382: T0 = 32'hf08f0006;
    383: T0 = 32'h59bf03d7;
    384: T0 = 32'h77bc3800;
    385: T0 = 32'h600302fb;
    386: T0 = 32'h8f1ff000;
    387: T0 = 32'h1e86d7fd;
    388: T0 = 32'h93c431b3;
    389: T0 = 32'h1f611e5d;
    390: T0 = 32'h7aac925f;
    391: T0 = 32'ha2207d19;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T5 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T6 = reset ? 1'h0 : restartRegs_0;
  assign T7 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_5(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T5;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T6;
  reg  restartRegs_0;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (addr)
    0: T0 = 32'ha4788037;
    1: T0 = 32'h7e2e66c3;
    2: T0 = 32'h1f634075;
    3: T0 = 32'hce5395e0;
    4: T0 = 32'h4f2f0017;
    5: T0 = 32'h8ecd89f5;
    6: T0 = 32'h304a000;
    7: T0 = 32'ha500000e;
    8: T0 = 32'h14b800;
    9: T0 = 32'hde000000;
    10: T0 = 32'h6010fd8;
    11: T0 = 32'hc4064f0;
    12: T0 = 32'h5b;
    13: T0 = 32'h5286fff;
    14: T0 = 32'hf200800d;
    15: T0 = 32'h32e249df;
    16: T0 = 32'h8ff8fb00;
    17: T0 = 32'hffff8073;
    18: T0 = 32'hf17f3fbe;
    19: T0 = 32'hfffffc87;
    20: T0 = 32'hf9ef3be3;
    21: T0 = 32'hff8f3fff;
    22: T0 = 32'hffc12458;
    23: T0 = 32'h69f023ff;
    24: T0 = 32'hafbcf667;
    25: T0 = 32'he9f81a1f;
    26: T0 = 32'h82ef7f3a;
    27: T0 = 32'hff579170;
    28: T0 = 32'h3fb703f9;
    29: T0 = 32'hfffb9587;
    30: T0 = 32'hb7f37817;
    31: T0 = 32'hfffe7810;
    32: T0 = 32'hdadf80c0;
    33: T0 = 32'hc8ff043b;
    34: T0 = 32'hf8bc98d0;
    35: T0 = 32'h94810045;
    36: T0 = 32'h611a9e0;
    37: T0 = 32'h3e000000;
    38: T0 = 32'haff;
    39: T0 = 32'h3b0f000;
    40: T0 = 32'hc0f053b7;
    41: T0 = 32'h21f1cb80;
    42: T0 = 32'hfc71030a;
    43: T0 = 32'h16d27e;
    44: T0 = 32'h55f20403;
    45: T0 = 32'hc806bd69;
    46: T0 = 32'h9017da04;
    47: T0 = 32'h9fee2887;
    48: T0 = 32'h67554c70;
    49: T0 = 32'hf2cf7c1f;
    50: T0 = 32'ha7930a;
    51: T0 = 32'h871e45d2;
    52: T0 = 32'ha084831a;
    53: T0 = 32'h4703682;
    54: T0 = 32'h79e902cb;
    55: T0 = 32'h8647d0cc;
    56: T0 = 32'h323cc121;
    57: T0 = 32'hf9fe2eff;
    58: T0 = 32'h89c0ff00;
    59: T0 = 32'h1f7e4127;
    60: T0 = 32'h7d08dbf8;
    61: T0 = 32'h93d0ef;
    62: T0 = 32'hf1b7edf;
    63: T0 = 32'hc000c5c4;
    64: T0 = 32'hc6fd37ef;
    65: T0 = 32'hb9031ea7;
    66: T0 = 32'h3e0fc37d;
    67: T0 = 32'hcc0c0f3;
    68: T0 = 32'h1f0f1e7;
    69: T0 = 32'he3c5fc07;
    70: T0 = 32'h260f7b6a;
    71: T0 = 32'h7a9fdfc0;
    72: T0 = 32'hdc4007ae;
    73: T0 = 32'h203686b0;
    74: T0 = 32'h63003a;
    75: T0 = 32'h7c0184e2;
    76: T0 = 32'hc62c003;
    77: T0 = 32'h87f43906;
    78: T0 = 32'hc1c45280;
    79: T0 = 32'he8fd0194;
    80: T0 = 32'h7c3d26c8;
    81: T0 = 32'h550fc002;
    82: T0 = 32'h79c1ff50;
    83: T0 = 32'h60a7c1;
    84: T0 = 32'hdcbcffe3;
    85: T0 = 32'he04396ff;
    86: T0 = 32'h1a0bffff;
    87: T0 = 32'hfe1bf87f;
    88: T0 = 32'h372fffe;
    89: T0 = 32'h17e0d3ac;
    90: T0 = 32'haaf7ff;
    91: T0 = 32'h807ffc0f;
    92: T0 = 32'hf80771df;
    93: T0 = 32'he4232000;
    94: T0 = 32'hffc1103c;
    95: T0 = 32'h1b17231c;
    96: T0 = 32'hdfff4e8e;
    97: T0 = 32'habeafa88;
    98: T0 = 32'h969833c2;
    99: T0 = 32'h21e181ed;
    100: T0 = 32'he75f6857;
    101: T0 = 32'h3b8ff001;
    102: T0 = 32'h917e3fe;
    103: T0 = 32'h57c5dbf3;
    104: T0 = 32'hf32d175f;
    105: T0 = 32'h4bff1fbb;
    106: T0 = 32'h270ced1b;
    107: T0 = 32'hbe000ff;
    108: T0 = 32'hfdd9b9da;
    109: T0 = 32'h80bef8ff;
    110: T0 = 32'h3fd4c03d;
    111: T0 = 32'h8953bebf;
    112: T0 = 32'hc4ac400f;
    113: T0 = 32'hc0102fb9;
    114: T0 = 32'h58010000;
    115: T0 = 32'h100000b8;
    116: T0 = 32'h22804000;
    117: T0 = 32'h220001c1;
    118: T0 = 32'hacbc1c;
    119: T0 = 32'h2230e040;
    120: T0 = 32'h301;
    121: T0 = 32'h5be4dfff;
    122: T0 = 32'h4000f197;
    123: T0 = 32'hf35e27ff;
    124: T0 = 32'hf000ffe8;
    125: T0 = 32'h3f73007f;
    126: T0 = 32'h6fc0fff6;
    127: T0 = 32'hff58803;
    128: T0 = 32'hc65e0fff;
    129: T0 = 32'hf1ffe480;
    130: T0 = 32'hfa2f0d7f;
    131: T0 = 32'heffffa14;
    132: T0 = 32'hffdf61d3;
    133: T0 = 32'h7eff0602;
    134: T0 = 32'hfff638f5;
    135: T0 = 32'h2bbff000;
    136: T0 = 32'hfbec0687;
    137: T0 = 32'hb38b840;
    138: T0 = 32'hffe0002c;
    139: T0 = 32'h26b0f84;
    140: T0 = 32'h57e07e0d;
    141: T0 = 32'h1253cafc;
    142: T0 = 32'h4cfef7f8;
    143: T0 = 32'h60b1b;
    144: T0 = 32'h5671fffb;
    145: T0 = 32'h38326351;
    146: T0 = 32'hbc2f4ede;
    147: T0 = 32'hc6c3b229;
    148: T0 = 32'h1ed85d83;
    149: T0 = 32'h776e40b3;
    150: T0 = 32'hdd3e2c4d;
    151: T0 = 32'he1a4200b;
    152: T0 = 32'he00e6f87;
    153: T0 = 32'hf4314400;
    154: T0 = 32'h7f838bcf;
    155: T0 = 32'h5eed2b5a;
    156: T0 = 32'hcf1e142f;
    157: T0 = 32'h61fcbb81;
    158: T0 = 32'h5d270001;
    159: T0 = 32'h3f070d4c;
    160: T0 = 32'h7f44d000;
    161: T0 = 32'h83f10054;
    162: T0 = 32'hff199fc;
    163: T0 = 32'h600ff807;
    164: T0 = 32'hf0fffb1f;
    165: T0 = 32'hf7c0ffff;
    166: T0 = 32'h7f87ffcd;
    167: T0 = 32'h3cf0cfff;
    168: T0 = 32'h2ff8fff8;
    169: T0 = 32'hc087ecff;
    170: T0 = 32'h45ff77ff;
    171: T0 = 32'hfe01f14b;
    172: T0 = 32'hefc01f;
    173: T0 = 32'hbbf87e11;
    174: T0 = 32'hc17e4e81;
    175: T0 = 32'h709f1932;
    176: T0 = 32'hbf8c88f8;
    177: T0 = 32'hdf0f80da;
    178: T0 = 32'h37fe0485;
    179: T0 = 32'hb0208d8f;
    180: T0 = 32'h8fff4280;
    181: T0 = 32'hf96e86a0;
    182: T0 = 32'hb48bc223;
    183: T0 = 32'h840ff90c;
    184: T0 = 32'he372ea88;
    185: T0 = 32'h10007711;
    186: T0 = 32'h2dd00f2b;
    187: T0 = 32'ha00ccff7;
    188: T0 = 32'he113ebd;
    189: T0 = 32'hde80ffe0;
    190: T0 = 32'h240545;
    191: T0 = 32'h60f8f27c;
    192: T0 = 32'h32004ea7;
    193: T0 = 32'h26e9ff76;
    194: T0 = 32'h17900ea6;
    195: T0 = 32'hf587d935;
    196: T0 = 32'hb7a06dc9;
    197: T0 = 32'h3b99ead3;
    198: T0 = 32'h690db050;
    199: T0 = 32'h3bd018e9;
    200: T0 = 32'heab6180c;
    201: T0 = 32'hac1e3e70;
    202: T0 = 32'heb3aa640;
    203: T0 = 32'h2037175c;
    204: T0 = 32'hffe7cc94;
    205: T0 = 32'h539f817f;
    206: T0 = 32'hfffeffef;
    207: T0 = 32'hdafffc07;
    208: T0 = 32'hffff17d1;
    209: T0 = 32'ha1fc183;
    210: T0 = 32'hafe039bb;
    211: T0 = 32'h298a7c;
    212: T0 = 32'h2000c3e5;
    213: T0 = 32'hf847;
    214: T0 = 32'h11817e0b;
    215: T0 = 32'h103f4;
    216: T0 = 32'h85487e0;
    217: T0 = 32'h100000d;
    218: T0 = 32'h1e41cc7f;
    219: T0 = 32'h49fef002;
    220: T0 = 32'hfffe18a3;
    221: T0 = 32'he00f1f80;
    222: T0 = 32'h2fff1840;
    223: T0 = 32'h2c36c1fc;
    224: T0 = 32'h3117e295;
    225: T0 = 32'h7f99727f;
    226: T0 = 32'h469efe01;
    227: T0 = 32'h55d93b7f;
    228: T0 = 32'h1a096fe0;
    229: T0 = 32'h998c0dc4;
    230: T0 = 32'h64a0d01c;
    231: T0 = 32'h63fec0d3;
    232: T0 = 32'hfdf73749;
    233: T0 = 32'h43fc023;
    234: T0 = 32'hffffb35f;
    235: T0 = 32'hfc973f82;
    236: T0 = 32'h7fff0db7;
    237: T0 = 32'hff4c7dd8;
    238: T0 = 32'h7bff01f2;
    239: T0 = 32'h5c2136f0;
    240: T0 = 32'he8ffc5f1;
    241: T0 = 32'h5e763;
    242: T0 = 32'h88c8b7cd;
    243: T0 = 32'h473e8236;
    244: T0 = 32'hfe6a4784;
    245: T0 = 32'h917b0c83;
    246: T0 = 32'h18d488c9;
    247: T0 = 32'h342fc045;
    248: T0 = 32'h8722c3f5;
    249: T0 = 32'h52f666bc;
    250: T0 = 32'hf013e007;
    251: T0 = 32'h7d863db;
    252: T0 = 32'hde000007;
    253: T0 = 32'h327abc81;
    254: T0 = 32'hf3e0f000;
    255: T0 = 32'h80c50690;
    256: T0 = 32'h5ffc816;
    257: T0 = 32'hfe734037;
    258: T0 = 32'hfc8f5f00;
    259: T0 = 32'hdfff0f85;
    260: T0 = 32'hfcc767f0;
    261: T0 = 32'h9fef01f8;
    262: T0 = 32'hf8018b7e;
    263: T0 = 32'h3ff403f;
    264: T0 = 32'hfd80fc5e;
    265: T0 = 32'hf78007;
    266: T0 = 32'hd778ffc7;
    267: T0 = 32'hfc072220;
    268: T0 = 32'h4c211ffc;
    269: T0 = 32'h3bfc0087;
    270: T0 = 32'he0a131f9;
    271: T0 = 32'h3f3fe1e0;
    272: T0 = 32'hfffc600f;
    273: T0 = 32'h41f1fe01;
    274: T0 = 32'hff9b000;
    275: T0 = 32'h827607f0;
    276: T0 = 32'h783f0fb0;
    277: T0 = 32'hfd17003f;
    278: T0 = 32'he003f8ef;
    279: T0 = 32'h1f1dc803;
    280: T0 = 32'h3c80ffc2;
    281: T0 = 32'h1f17500;
    282: T0 = 32'hcde8fe30;
    283: T0 = 32'h801ef8fb;
    284: T0 = 32'he56cffbf;
    285: T0 = 32'hcc031da2;
    286: T0 = 32'hfcf2aff9;
    287: T0 = 32'h7b001b5c;
    288: T0 = 32'h7f044b7f;
    289: T0 = 32'hc4f75243;
    290: T0 = 32'h9fe0d58e;
    291: T0 = 32'h899ba102;
    292: T0 = 32'h4bc053ce;
    293: T0 = 32'h122e28a1;
    294: T0 = 32'hecb291ad;
    295: T0 = 32'hddc09df2;
    296: T0 = 32'hb381dd64;
    297: T0 = 32'hf0c13647;
    298: T0 = 32'h488ed29f;
    299: T0 = 32'h30653a0f;
    300: T0 = 32'he44cc200;
    301: T0 = 32'h7e1fff3d;
    302: T0 = 32'hdff15189;
    303: T0 = 32'h48fb7f24;
    304: T0 = 32'hcdfb0f0e;
    305: T0 = 32'hfbba5ffe;
    306: T0 = 32'h6cfff0f5;
    307: T0 = 32'hfeb487ff;
    308: T0 = 32'h786ff8d;
    309: T0 = 32'he7e8fccf;
    310: T0 = 32'hc4a07fe;
    311: T0 = 32'h387ff374;
    312: T0 = 32'hff80000f;
    313: T0 = 32'h387073e;
    314: T0 = 32'h7fd0b2dc;
    315: T0 = 32'h140c03f;
    316: T0 = 32'h7f2cbff;
    317: T0 = 32'h563cce00;
    318: T0 = 32'he07e0ef9;
    319: T0 = 32'hc68700f0;
    320: T0 = 32'hcfc70117;
    321: T0 = 32'hf871100f;
    322: T0 = 32'h9fd6fc3a;
    323: T0 = 32'h7f863883;
    324: T0 = 32'h79f10f27;
    325: T0 = 32'hff1f4da;
    326: T0 = 32'h121fb064;
    327: T0 = 32'hf87c1ffd;
    328: T0 = 32'h4cfe06;
    329: T0 = 32'hcf8103ef;
    330: T0 = 32'h3003b73a;
    331: T0 = 32'h2afc80ff;
    332: T0 = 32'he030a87f;
    333: T0 = 32'hb68fe65f;
    334: T0 = 32'hff01100b;
    335: T0 = 32'h624153a;
    336: T0 = 32'hebf8fa26;
    337: T0 = 32'heaca763f;
    338: T0 = 32'h3d5ffffd;
    339: T0 = 32'hfffe0255;
    340: T0 = 32'hc68f7ff4;
    341: T0 = 32'h767f6cf7;
    342: T0 = 32'h79ed01c4;
    343: T0 = 32'h372600bc;
    344: T0 = 32'hafe5ba8;
    345: T0 = 32'ha515b04;
    346: T0 = 32'hb7f679a2;
    347: T0 = 32'hfbd1fe02;
    348: T0 = 32'hbd0e376a;
    349: T0 = 32'h3ea789c0;
    350: T0 = 32'hbc000a53;
    351: T0 = 32'h1fc1e55e;
    352: T0 = 32'h8fab01ae;
    353: T0 = 32'hf1e0fbce;
    354: T0 = 32'h1480f03f;
    355: T0 = 32'h2718f963;
    356: T0 = 32'h1bde7dc3;
    357: T0 = 32'hacf83ffc;
    358: T0 = 32'h6fa2ffc;
    359: T0 = 32'hfc77c1fb;
    360: T0 = 32'hf83feb7f;
    361: T0 = 32'hfec2fc3c;
    362: T0 = 32'hff87ffd7;
    363: T0 = 32'h3dc4af6f;
    364: T0 = 32'h9ffcfff7;
    365: T0 = 32'he0aa7605;
    366: T0 = 32'h15ffbfff;
    367: T0 = 32'h7f808900;
    368: T0 = 32'h17f2fff;
    369: T0 = 32'hfbf88034;
    370: T0 = 32'hc257047f;
    371: T0 = 32'h5e9ff006;
    372: T0 = 32'h7ded6803;
    373: T0 = 32'hb70e00;
    374: T0 = 32'hffff0700;
    375: T0 = 32'hf4051000;
    376: T0 = 32'h7ff0060;
    377: T0 = 32'hff4cc000;
    378: T0 = 32'hf03f0005;
    379: T0 = 32'h1ff24800;
    380: T0 = 32'hd500000b;
    381: T0 = 32'hb7780;
    382: T0 = 32'hb10038d6;
    383: T0 = 32'h1800ac20;
    384: T0 = 32'h839840ff;
    385: T0 = 32'hca80ff18;
    386: T0 = 32'h202f4637;
    387: T0 = 32'he09fff6;
    388: T0 = 32'h415e7;
    389: T0 = 32'h93409fa0;
    390: T0 = 32'he4003637;
    391: T0 = 32'h4c126377;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T5 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T6 = reset ? 1'h0 : restartRegs_0;
  assign T7 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_6(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T5;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T6;
  reg  restartRegs_0;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (addr)
    0: T0 = 32'h2f455842;
    1: T0 = 32'hb814643b;
    2: T0 = 32'h6ccff05b;
    3: T0 = 32'h684139d0;
    4: T0 = 32'h8d51eecb;
    5: T0 = 32'h20611174;
    6: T0 = 32'h11c1f64;
    7: T0 = 32'h8009fdc;
    8: T0 = 32'h7829fe;
    9: T0 = 32'h9b0fe0a;
    10: T0 = 32'h80017ac1;
    11: T0 = 32'h119f0098;
    12: T0 = 32'hffc06fbc;
    13: T0 = 32'h8041fc00;
    14: T0 = 32'h1fff01e2;
    15: T0 = 32'hfd8053f8;
    16: T0 = 32'h77fff91;
    17: T0 = 32'h7fbe10ff;
    18: T0 = 32'hf0807ffd;
    19: T0 = 32'hfff673;
    20: T0 = 32'hff2c81ff;
    21: T0 = 32'hc00cff9f;
    22: T0 = 32'hc3f2580f;
    23: T0 = 32'hfe3c7f91;
    24: T0 = 32'hfc3f22a0;
    25: T0 = 32'h1ea103f0;
    26: T0 = 32'he000ac;
    27: T0 = 32'he44a9e;
    28: T0 = 32'h8006801a;
    29: T0 = 32'h7000b7e8;
    30: T0 = 32'h82007803;
    31: T0 = 32'hf84da8d;
    32: T0 = 32'h8e806b80;
    33: T0 = 32'h4fc07a8;
    34: T0 = 32'he00e8378;
    35: T0 = 32'h70dec35b;
    36: T0 = 32'h4328381f;
    37: T0 = 32'he0f7820;
    38: T0 = 32'h804247e0;
    39: T0 = 32'hf15f0f88;
    40: T0 = 32'hff418b05;
    41: T0 = 32'h873fe0fd;
    42: T0 = 32'h3fd0cfd1;
    43: T0 = 32'hdb89530f;
    44: T0 = 32'h6e7f7ffc;
    45: T0 = 32'hfffe1368;
    46: T0 = 32'hd8fac7eb;
    47: T0 = 32'hf3ffd176;
    48: T0 = 32'h82222ab5;
    49: T0 = 32'h16b081f9;
    50: T0 = 32'hb907e464;
    51: T0 = 32'h2e0946cb;
    52: T0 = 32'h10fcb44d;
    53: T0 = 32'h92d0e5c;
    54: T0 = 32'h9b835cf2;
    55: T0 = 32'h10a9f838;
    56: T0 = 32'h89b0e611;
    57: T0 = 32'h198600;
    58: T0 = 32'h79fd0f1e;
    59: T0 = 32'h8000a318;
    60: T0 = 32'h1dfc0eb;
    61: T0 = 32'h78f0035f;
    62: T0 = 32'hc0723f0e;
    63: T0 = 32'h6f8fe23e;
    64: T0 = 32'h7f1e77ff;
    65: T0 = 32'h76b8fe05;
    66: T0 = 32'hc3f88b5f;
    67: T0 = 32'h9ec7fff0;
    68: T0 = 32'h7e0f009f;
    69: T0 = 32'h5fc61fcf;
    70: T0 = 32'h17f0f007;
    71: T0 = 32'h807d4b80;
    72: T0 = 32'hd4ff0f80;
    73: T0 = 32'hfc0102b8;
    74: T0 = 32'h288700fc;
    75: T0 = 32'h3ff9973b;
    76: T0 = 32'h83ec810f;
    77: T0 = 32'hdfffe12;
    78: T0 = 32'hfdbc9880;
    79: T0 = 32'hd9c3075c;
    80: T0 = 32'h1fd3f16d;
    81: T0 = 32'h1edcc87d;
    82: T0 = 32'he8de78;
    83: T0 = 32'h3651df67;
    84: T0 = 32'h18003fc8;
    85: T0 = 32'hf0c868;
    86: T0 = 32'he40023f9;
    87: T0 = 32'h963ce66;
    88: T0 = 32'hf788481f;
    89: T0 = 32'h10ff8a;
    90: T0 = 32'h22c0a8;
    91: T0 = 32'h14034fc6;
    92: T0 = 32'he30a6340;
    93: T0 = 32'hdc0008bf;
    94: T0 = 32'hfffed962;
    95: T0 = 32'h8f183f98;
    96: T0 = 32'h97895acf;
    97: T0 = 32'h797ea5dc;
    98: T0 = 32'hd8677efa;
    99: T0 = 32'h97f7ead1;
    100: T0 = 32'h8fc1cd42;
    101: T0 = 32'hdc3759dc;
    102: T0 = 32'h4de4d7fd;
    103: T0 = 32'hf80dbb06;
    104: T0 = 32'h473609de;
    105: T0 = 32'hebd9264f;
    106: T0 = 32'hbdcc76;
    107: T0 = 32'h941ee201;
    108: T0 = 32'hf5224bf6;
    109: T0 = 32'h11542f20;
    110: T0 = 32'h898e8580;
    111: T0 = 32'hb438643;
    112: T0 = 32'h80000028;
    113: T0 = 32'ha69453;
    114: T0 = 32'hbc00f140;
    115: T0 = 32'hff0185;
    116: T0 = 32'hfc401e01;
    117: T0 = 32'he07f0070;
    118: T0 = 32'hff0d0fc0;
    119: T0 = 32'h3fdf080b;
    120: T0 = 32'hfff491e8;
    121: T0 = 32'ha6ff801e;
    122: T0 = 32'hffbff8be;
    123: T0 = 32'hf2bff807;
    124: T0 = 32'hfff9ff29;
    125: T0 = 32'h80977fc0;
    126: T0 = 32'hffff3ff1;
    127: T0 = 32'hfd0937fe;
    128: T0 = 32'h3ffbe3fe;
    129: T0 = 32'h7e08627;
    130: T0 = 32'h7be7f1f;
    131: T0 = 32'h7ee42b;
    132: T0 = 32'h7541f1;
    133: T0 = 32'he0008f2a;
    134: T0 = 32'h48b93;
    135: T0 = 32'h3400f8f8;
    136: T0 = 32'h1440bd3f;
    137: T0 = 32'had22f703;
    138: T0 = 32'h892c3edd;
    139: T0 = 32'h9e15bc60;
    140: T0 = 32'hf22103ac;
    141: T0 = 32'he29ff8f;
    142: T0 = 32'h180dd01f;
    143: T0 = 32'h8202f356;
    144: T0 = 32'h12ccd889;
    145: T0 = 32'h2808b1f0;
    146: T0 = 32'ha164bf4c;
    147: T0 = 32'h8f45811d;
    148: T0 = 32'h95d3d6ab;
    149: T0 = 32'h7580e172;
    150: T0 = 32'h28d13513;
    151: T0 = 32'hebb7712a;
    152: T0 = 32'h60fd8726;
    153: T0 = 32'h2dc19f8e;
    154: T0 = 32'h4cc1137b;
    155: T0 = 32'h1fc5f6f8;
    156: T0 = 32'h13f0a0fe;
    157: T0 = 32'h7fe00f;
    158: T0 = 32'hfe3fbf87;
    159: T0 = 32'hd07f3f9f;
    160: T0 = 32'hff37b5fc;
    161: T0 = 32'hdd07c3f7;
    162: T0 = 32'h1fffc41f;
    163: T0 = 32'h5f503c3f;
    164: T0 = 32'h384e6200;
    165: T0 = 32'h647a01c3;
    166: T0 = 32'h3c17e2a;
    167: T0 = 32'h8107403c;
    168: T0 = 32'h607fc7fa;
    169: T0 = 32'hff07ea07;
    170: T0 = 32'h9007dc3b;
    171: T0 = 32'h35ff7f80;
    172: T0 = 32'h21401fc0;
    173: T0 = 32'hb010b38;
    174: T0 = 32'h49866ec;
    175: T0 = 32'h407c40ca;
    176: T0 = 32'h701fa291;
    177: T0 = 32'hc0162601;
    178: T0 = 32'hf7031910;
    179: T0 = 32'h36801ee0;
    180: T0 = 32'h17380710;
    181: T0 = 32'h8294a27f;
    182: T0 = 32'he1f7f032;
    183: T0 = 32'h781c7807;
    184: T0 = 32'h863fff01;
    185: T0 = 32'hbb891518;
    186: T0 = 32'hcbfefe1;
    187: T0 = 32'hf3f03ee9;
    188: T0 = 32'h2fe4eff8;
    189: T0 = 32'h57fc01f7;
    190: T0 = 32'hc2fb70ff;
    191: T0 = 32'h2c7f4aff;
    192: T0 = 32'hf806dc62;
    193: T0 = 32'h4c5ff6df;
    194: T0 = 32'hcc02a91c;
    195: T0 = 32'h218a8f10;
    196: T0 = 32'hd64c35b1;
    197: T0 = 32'h9f201b17;
    198: T0 = 32'hea6e2cfb;
    199: T0 = 32'h67dcb8c;
    200: T0 = 32'h7ed6dc0;
    201: T0 = 32'h445a001f;
    202: T0 = 32'hc9c67260;
    203: T0 = 32'h6c07c028;
    204: T0 = 32'h7f674c5f;
    205: T0 = 32'h1180b700;
    206: T0 = 32'h1bde4f3;
    207: T0 = 32'h42d0be37;
    208: T0 = 32'h1fffec;
    209: T0 = 32'h2f4607fb;
    210: T0 = 32'h601c3ffe;
    211: T0 = 32'hf4bf6aff;
    212: T0 = 32'ha203f078;
    213: T0 = 32'h3f4b01cd;
    214: T0 = 32'hb9401f00;
    215: T0 = 32'h1f44028;
    216: T0 = 32'h3d917f8;
    217: T0 = 32'h840fc00e;
    218: T0 = 32'h611ca63f;
    219: T0 = 32'hea0ff01;
    220: T0 = 32'hc0031e83;
    221: T0 = 32'h18af0ff8;
    222: T0 = 32'hfe00f7f6;
    223: T0 = 32'h28f620ff;
    224: T0 = 32'hf7f8fffd;
    225: T0 = 32'hc086d883;
    226: T0 = 32'h37fd3fff;
    227: T0 = 32'hfe08f688;
    228: T0 = 32'h5b7f103f;
    229: T0 = 32'hfbe06590;
    230: T0 = 32'h4f4300;
    231: T0 = 32'hbfa6001e;
    232: T0 = 32'h7000c8d0;
    233: T0 = 32'hd6c00007;
    234: T0 = 32'h2b00dc5a;
    235: T0 = 32'h920ff41;
    236: T0 = 32'h82dc0412;
    237: T0 = 32'hc05db7f2;
    238: T0 = 32'h703f2816;
    239: T0 = 32'hfc0c4938;
    240: T0 = 32'ha5b0841;
    241: T0 = 32'h7ff09c69;
    242: T0 = 32'h87848805;
    243: T0 = 32'hcfcf175c;
    244: T0 = 32'h8aba4037;
    245: T0 = 32'hf406aeff;
    246: T0 = 32'h356981f0;
    247: T0 = 32'h3cba8087;
    248: T0 = 32'hc19b7bd4;
    249: T0 = 32'hf3cb1789;
    250: T0 = 32'h9e6fa8ca;
    251: T0 = 32'hdc1ad07f;
    252: T0 = 32'h8113fe78;
    253: T0 = 32'h37ee7f41;
    254: T0 = 32'hc205deb;
    255: T0 = 32'h23783c4;
    256: T0 = 32'h7d605fff;
    257: T0 = 32'hb4e2d0;
    258: T0 = 32'h3facaff;
    259: T0 = 32'h4000fc49;
    260: T0 = 32'h3e23203;
    261: T0 = 32'hdb300140;
    262: T0 = 32'hfc150fa0;
    263: T0 = 32'h6bf4000;
    264: T0 = 32'hffe080aa;
    265: T0 = 32'h8b87bff1;
    266: T0 = 32'hbffffd5a;
    267: T0 = 32'hfc2543ff;
    268: T0 = 32'heffffffe;
    269: T0 = 32'hffc8faff;
    270: T0 = 32'h631dffbf;
    271: T0 = 32'hfffeff13;
    272: T0 = 32'hfd6b7ff9;
    273: T0 = 32'h7fff0ff4;
    274: T0 = 32'hfde04fff;
    275: T0 = 32'he5ff807f;
    276: T0 = 32'hffeffc7f;
    277: T0 = 32'hf29ff603;
    278: T0 = 32'h7fff1eab;
    279: T0 = 32'hfd88fe00;
    280: T0 = 32'h109f0076;
    281: T0 = 32'h59eec00;
    282: T0 = 32'h71000008;
    283: T0 = 32'h40abe;
    284: T0 = 32'ha390e086;
    285: T0 = 32'h209811;
    286: T0 = 32'h104e6800;
    287: T0 = 32'he04f05f4;
    288: T0 = 32'h127640;
    289: T0 = 32'h6815be2f;
    290: T0 = 32'h44c359d;
    291: T0 = 32'h82b20ff4;
    292: T0 = 32'he8029d16;
    293: T0 = 32'h9d900fc7;
    294: T0 = 32'hcc800614;
    295: T0 = 32'hbe8fa79e;
    296: T0 = 32'h6371581;
    297: T0 = 32'hc7b7836e;
    298: T0 = 32'h3100402a;
    299: T0 = 32'he806734d;
    300: T0 = 32'h293cffe5;
    301: T0 = 32'h4580bf1a;
    302: T0 = 32'h106d734;
    303: T0 = 32'h34fcfff6;
    304: T0 = 32'h8001c2c3;
    305: T0 = 32'h189dffff;
    306: T0 = 32'he01cfe6e;
    307: T0 = 32'hfd1dd403;
    308: T0 = 32'hfe010f61;
    309: T0 = 32'h3fff2420;
    310: T0 = 32'hbbc0001b;
    311: T0 = 32'h7ff0159;
    312: T0 = 32'hfa784001;
    313: T0 = 32'h807f4a70;
    314: T0 = 32'hffef1900;
    315: T0 = 32'h3c071d43;
    316: T0 = 32'hf9fc55ff;
    317: T0 = 32'h43c0f9e0;
    318: T0 = 32'hfcf847f;
    319: T0 = 32'h107effbd;
    320: T0 = 32'hf07ec06b;
    321: T0 = 32'h39b71fff;
    322: T0 = 32'hff87ffc5;
    323: T0 = 32'he3c0b5ff;
    324: T0 = 32'hf7fcfff2;
    325: T0 = 32'he6dcfd1f;
    326: T0 = 32'he67f7d9e;
    327: T0 = 32'h72808fc3;
    328: T0 = 32'h682aff8;
    329: T0 = 32'h200e90f8;
    330: T0 = 32'hb263016e;
    331: T0 = 32'h7204ffff;
    332: T0 = 32'h88c8e2e3;
    333: T0 = 32'ha6a01dff;
    334: T0 = 32'hdf10c13e;
    335: T0 = 32'h387c1eff;
    336: T0 = 32'h2af8ff39;
    337: T0 = 32'h2926bfc;
    338: T0 = 32'h37e0041;
    339: T0 = 32'he003c2e4;
    340: T0 = 32'h4067c00c;
    341: T0 = 32'h7e00d2c9;
    342: T0 = 32'h398e4a20;
    343: T0 = 32'hf84316d;
    344: T0 = 32'h9ffac0ba;
    345: T0 = 32'hbc740913;
    346: T0 = 32'h8c95e0d6;
    347: T0 = 32'h209fec12;
    348: T0 = 32'h400740dc;
    349: T0 = 32'hd7373b40;
    350: T0 = 32'he06d0058;
    351: T0 = 32'h8af395ef;
    352: T0 = 32'hd447000;
    353: T0 = 32'h270162cf;
    354: T0 = 32'ha1cfc1f;
    355: T0 = 32'h3ffcff9f;
    356: T0 = 32'hf0987fc0;
    357: T0 = 32'h93ff1ffc;
    358: T0 = 32'hffd49be0;
    359: T0 = 32'h6d1503ff;
    360: T0 = 32'h3fd97bb8;
    361: T0 = 32'h23c0003f;
    362: T0 = 32'h77fef3f2;
    363: T0 = 32'h9ed86003;
    364: T0 = 32'hafff1d98;
    365: T0 = 32'hf06dc600;
    366: T0 = 32'hedff00e6;
    367: T0 = 32'hf0039740;
    368: T0 = 32'h37f5c05;
    369: T0 = 32'hfe002c24;
    370: T0 = 32'h37ff8;
    371: T0 = 32'hbfe0c08c;
    372: T0 = 32'h1433f;
    373: T0 = 32'h2bfffc0e;
    374: T0 = 32'hf038f47b;
    375: T0 = 32'h155ff7e0;
    376: T0 = 32'h76050f9f;
    377: T0 = 32'h5fcffe0e;
    378: T0 = 32'h80e0ff;
    379: T0 = 32'h3ffc5e1;
    380: T0 = 32'hf808b8c1;
    381: T0 = 32'hfd1fe;
    382: T0 = 32'h8e70ff9e;
    383: T0 = 32'h19515b;
    384: T0 = 32'hff049e3c;
    385: T0 = 32'h900f7a54;
    386: T0 = 32'h3ff25900;
    387: T0 = 32'h7c800100;
    388: T0 = 32'hfffe0c88;
    389: T0 = 32'hee27d38e;
    390: T0 = 32'h6263391f;
    391: T0 = 32'h909f3560;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T5 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T6 = reset ? 1'h0 : restartRegs_0;
  assign T7 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_7(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T5;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T6;
  reg  restartRegs_0;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (addr)
    0: T0 = 32'h232927c5;
    1: T0 = 32'hf7043146;
    2: T0 = 32'hebbad895;
    3: T0 = 32'h83915bc7;
    4: T0 = 32'h2fea9a90;
    5: T0 = 32'h76694;
    6: T0 = 32'hd666cdc0;
    7: T0 = 32'h501e013b;
    8: T0 = 32'h7e63fed3;
    9: T0 = 32'h3e04e00f;
    10: T0 = 32'hffc0654e;
    11: T0 = 32'h726f800;
    12: T0 = 32'hf7f03156;
    13: T0 = 32'h9ea000;
    14: T0 = 32'hcff3ff3;
    15: T0 = 32'hc013f040;
    16: T0 = 32'h46ff07ff;
    17: T0 = 32'hf801fa00;
    18: T0 = 32'hb4f00ff;
    19: T0 = 32'hff00feb0;
    20: T0 = 32'h1a78c1f;
    21: T0 = 32'hb9e0ffb3;
    22: T0 = 32'h32c9ef;
    23: T0 = 32'h945c3f04;
    24: T0 = 32'hc001eaff;
    25: T0 = 32'hf8aaf9fb;
    26: T0 = 32'h9c00fe07;
    27: T0 = 32'h3fa9ffaf;
    28: T0 = 32'hd3c0ffc7;
    29: T0 = 32'h7fd65ff;
    30: T0 = 32'he416fff8;
    31: T0 = 32'he1ff063f;
    32: T0 = 32'hfb10b25f;
    33: T0 = 32'hff3f006c;
    34: T0 = 32'hff3c7000;
    35: T0 = 32'h3fffc00a;
    36: T0 = 32'h9b712218;
    37: T0 = 32'h27eb4f49;
    38: T0 = 32'hfe44c320;
    39: T0 = 32'h843e0314;
    40: T0 = 32'hfff37d35;
    41: T0 = 32'hc1a1903f;
    42: T0 = 32'h9ffdff96;
    43: T0 = 32'hf75c1;
    44: T0 = 32'h98ffdfc8;
    45: T0 = 32'he000a5dd;
    46: T0 = 32'h96dbb980;
    47: T0 = 32'h7400cc2c;
    48: T0 = 32'h19ef3202;
    49: T0 = 32'h83997a4e;
    50: T0 = 32'h3ac7d9b1;
    51: T0 = 32'he9744c17;
    52: T0 = 32'hd9d1043a;
    53: T0 = 32'hef19ddd8;
    54: T0 = 32'h50339890;
    55: T0 = 32'h484f753f;
    56: T0 = 32'h40ffffe0;
    57: T0 = 32'he0d9567b;
    58: T0 = 32'h2e1f7ff7;
    59: T0 = 32'hf84927c1;
    60: T0 = 32'hb7c31fe1;
    61: T0 = 32'h7e0100f0;
    62: T0 = 32'h401603fc;
    63: T0 = 32'h6fe08000;
    64: T0 = 32'h183b05f;
    65: T0 = 32'hdf8f800;
    66: T0 = 32'h10090f;
    67: T0 = 32'h431fff00;
    68: T0 = 32'hf00e002c;
    69: T0 = 32'hff67cfe0;
    70: T0 = 32'h7f030408;
    71: T0 = 32'h3ff658fa;
    72: T0 = 32'hf7f0e07e;
    73: T0 = 32'h81ffebcf;
    74: T0 = 32'hf9cfb603;
    75: T0 = 32'hf89f9f08;
    76: T0 = 32'hfff041b0;
    77: T0 = 32'h1fe10374;
    78: T0 = 32'h81fa9803;
    79: T0 = 32'h841f9059;
    80: T0 = 32'h3e1ffe00;
    81: T0 = 32'hf2010045;
    82: T0 = 32'ha3e19f50;
    83: T0 = 32'h1f74c003;
    84: T0 = 32'hc2effb18;
    85: T0 = 32'hb1f5ca01;
    86: T0 = 32'hbae5fb87;
    87: T0 = 32'h67bfe6d7;
    88: T0 = 32'h78f56fdf;
    89: T0 = 32'he7becbb0;
    90: T0 = 32'h5839957f;
    91: T0 = 32'he0a0fdfe;
    92: T0 = 32'hcbdb59eb;
    93: T0 = 32'h1e1907df;
    94: T0 = 32'hbcffa2ac;
    95: T0 = 32'he864816f;
    96: T0 = 32'h3149dda1;
    97: T0 = 32'h7ae6868f;
    98: T0 = 32'h49265f1;
    99: T0 = 32'h91cedfa3;
    100: T0 = 32'h136988b2;
    101: T0 = 32'hb903f1dd;
    102: T0 = 32'hd8d500fd;
    103: T0 = 32'h185ca9b6;
    104: T0 = 32'he8edabff;
    105: T0 = 32'hc080c0c8;
    106: T0 = 32'hf95523f;
    107: T0 = 32'h599af801;
    108: T0 = 32'h8600219f;
    109: T0 = 32'h41cfed0;
    110: T0 = 32'h8070d245;
    111: T0 = 32'h81adefc0;
    112: T0 = 32'h9c0301c5;
    113: T0 = 32'h780667fc;
    114: T0 = 32'hfc0c0fa;
    115: T0 = 32'h380ea3f;
    116: T0 = 32'h3fdefc0f;
    117: T0 = 32'h54383fff;
    118: T0 = 32'h80b3ff80;
    119: T0 = 32'hbcc130f8;
    120: T0 = 32'h38061c78;
    121: T0 = 32'hbfc0830f;
    122: T0 = 32'h3c0fdc7;
    123: T0 = 32'h84fc7874;
    124: T0 = 32'hc23f0fc4;
    125: T0 = 32'hf679c3c3;
    126: T0 = 32'h9ea30cfc;
    127: T0 = 32'hbff8781c;
    128: T0 = 32'hfbdfe1ef;
    129: T0 = 32'hf9ffbee0;
    130: T0 = 32'hf83d0f9f;
    131: T0 = 32'hffdffe90;
    132: T0 = 32'hffc580fd;
    133: T0 = 32'h7fffeffe;
    134: T0 = 32'hdf7eb03e;
    135: T0 = 32'hcf3ffe3f;
    136: T0 = 32'h3bffb4f;
    137: T0 = 32'hffa2ff75;
    138: T0 = 32'h1f4e13;
    139: T0 = 32'he9a0cfdc;
    140: T0 = 32'hfe19;
    141: T0 = 32'h1e82fd;
    142: T0 = 32'h2400dfe1;
    143: T0 = 32'h4ca9f;
    144: T0 = 32'hbccf06f;
    145: T0 = 32'h9ff48766;
    146: T0 = 32'hf159e7fe;
    147: T0 = 32'ha9998767;
    148: T0 = 32'h5dd947f6;
    149: T0 = 32'hfa7f4996;
    150: T0 = 32'hd4453e5b;
    151: T0 = 32'hc5b2fef3;
    152: T0 = 32'h603dfd6e;
    153: T0 = 32'hfa68dfbf;
    154: T0 = 32'h1d01ff2a;
    155: T0 = 32'hb736eb7;
    156: T0 = 32'h22ecfffe;
    157: T0 = 32'h203ff787;
    158: T0 = 32'hf879ef99;
    159: T0 = 32'hc00f0fb7;
    160: T0 = 32'hfad10000;
    161: T0 = 32'hdff0003f;
    162: T0 = 32'h76fec00;
    163: T0 = 32'hc2ff0401;
    164: T0 = 32'hf8771880;
    165: T0 = 32'hfffbc3ff;
    166: T0 = 32'hffcfe4a5;
    167: T0 = 32'hff19ffef;
    168: T0 = 32'hfe78fc8d;
    169: T0 = 32'hff4fffe;
    170: T0 = 32'h87f08602;
    171: T0 = 32'hff033f;
    172: T0 = 32'hfd8ef800;
    173: T0 = 32'hda07064f;
    174: T0 = 32'h7b546f04;
    175: T0 = 32'h2400402;
    176: T0 = 32'h7495dc0;
    177: T0 = 32'h2c0001e6;
    178: T0 = 32'h2072e3a0;
    179: T0 = 32'h341913f;
    180: T0 = 32'h1fffda;
    181: T0 = 32'hc820af7f;
    182: T0 = 32'h8141ffe8;
    183: T0 = 32'h3c06245f;
    184: T0 = 32'h58087fff;
    185: T0 = 32'h1e8e9b2;
    186: T0 = 32'h66349fef;
    187: T0 = 32'hc81ef07f;
    188: T0 = 32'hfa50f47f;
    189: T0 = 32'h1c036213;
    190: T0 = 32'h7e0b6000;
    191: T0 = 32'h8f288000;
    192: T0 = 32'ha7038498;
    193: T0 = 32'h44f1abc6;
    194: T0 = 32'hc4e09167;
    195: T0 = 32'hf7a55341;
    196: T0 = 32'hfa71c7cb;
    197: T0 = 32'hafcf3dd4;
    198: T0 = 32'h6a62639c;
    199: T0 = 32'hd8e0bafc;
    200: T0 = 32'h59dba9ff;
    201: T0 = 32'h6ffdecb5;
    202: T0 = 32'hfbbaae07;
    203: T0 = 32'hafff2fd5;
    204: T0 = 32'hffe563c0;
    205: T0 = 32'h6be683f5;
    206: T0 = 32'h53fc761f;
    207: T0 = 32'hf4b0fc1d;
    208: T0 = 32'hffffc7a6;
    209: T0 = 32'h2e9f8c81;
    210: T0 = 32'h75ff0ffc;
    211: T0 = 32'h82bf808c;
    212: T0 = 32'h1811e1cf;
    213: T0 = 32'h2780b;
    214: T0 = 32'h1f80de1c;
    215: T0 = 32'h4000e750;
    216: T0 = 32'he60fe1;
    217: T0 = 32'h28000fce;
    218: T0 = 32'h381b5fe7;
    219: T0 = 32'h58e0707f;
    220: T0 = 32'h3f7f7bf;
    221: T0 = 32'he87fc303;
    222: T0 = 32'hf01f3bcf;
    223: T0 = 32'hfabbff20;
    224: T0 = 32'h3fc081dc;
    225: T0 = 32'he553e0;
    226: T0 = 32'h3ffc6c1e;
    227: T0 = 32'hf00bd6fe;
    228: T0 = 32'h17af7f61;
    229: T0 = 32'hff800e62;
    230: T0 = 32'hf3c280a4;
    231: T0 = 32'hfffb225;
    232: T0 = 32'hfffdae0e;
    233: T0 = 32'h467fa8e2;
    234: T0 = 32'h3fffcf21;
    235: T0 = 32'hfaa22827;
    236: T0 = 32'h803f3e52;
    237: T0 = 32'h3f201002;
    238: T0 = 32'h500087c1;
    239: T0 = 32'hdff9a202;
    240: T0 = 32'h7435276f;
    241: T0 = 32'he00b01e8;
    242: T0 = 32'hfa54cf86;
    243: T0 = 32'hbd30f6cf;
    244: T0 = 32'hceb4cb48;
    245: T0 = 32'h4fc9bd70;
    246: T0 = 32'h5f2519cf;
    247: T0 = 32'hac16dcba;
    248: T0 = 32'h489d6fdd;
    249: T0 = 32'hfda6daf4;
    250: T0 = 32'h4540fae6;
    251: T0 = 32'h558555f;
    252: T0 = 32'h40783e1a;
    253: T0 = 32'hf8053380;
    254: T0 = 32'hd40f0350;
    255: T0 = 32'hfffa8e7e;
    256: T0 = 32'hdac3d07f;
    257: T0 = 32'h3e07f80b;
    258: T0 = 32'h1d743907;
    259: T0 = 32'h3c07b6f;
    260: T0 = 32'hff3eff0;
    261: T0 = 32'h981c07de;
    262: T0 = 32'hf001eb3e;
    263: T0 = 32'h168080ff;
    264: T0 = 32'hf80f6c7;
    265: T0 = 32'hd4019f;
    266: T0 = 32'h807cff7c;
    267: T0 = 32'hd00e203f;
    268: T0 = 32'h1a01fff1;
    269: T0 = 32'h6f000183;
    270: T0 = 32'h11b507fc;
    271: T0 = 32'hfff80020;
    272: T0 = 32'h3fd3001f;
    273: T0 = 32'h5fdfc000;
    274: T0 = 32'hf3fb0c01;
    275: T0 = 32'hfbff0c00;
    276: T0 = 32'hff1b6e18;
    277: T0 = 32'h7c7f40e0;
    278: T0 = 32'h33e00fc0;
    279: T0 = 32'h798d99e;
    280: T0 = 32'hc000e097;
    281: T0 = 32'h7c7e41;
    282: T0 = 32'h70003e10;
    283: T0 = 32'hfc04876a;
    284: T0 = 32'h94a381e1;
    285: T0 = 32'h3ff80261;
    286: T0 = 32'h8ab98cbc;
    287: T0 = 32'h79ffc3c9;
    288: T0 = 32'hf152e353;
    289: T0 = 32'hc301fffe;
    290: T0 = 32'h1fe4e3;
    291: T0 = 32'h51f04fdb;
    292: T0 = 32'h40070735;
    293: T0 = 32'he3b5e0e7;
    294: T0 = 32'he334fce9;
    295: T0 = 32'h9956ddf4;
    296: T0 = 32'h5a5d8676;
    297: T0 = 32'hae1ba0a0;
    298: T0 = 32'h3a7157d0;
    299: T0 = 32'h24df0752;
    300: T0 = 32'ha2f3ddfd;
    301: T0 = 32'h6ccb08ff;
    302: T0 = 32'hf2cb30ff;
    303: T0 = 32'h9d8260aa;
    304: T0 = 32'h9f1c053f;
    305: T0 = 32'hf6b1ff83;
    306: T0 = 32'h1e3fa61;
    307: T0 = 32'h1fc51fa1;
    308: T0 = 32'h503e3fac;
    309: T0 = 32'he3d0fff0;
    310: T0 = 32'h76101fc;
    311: T0 = 32'hbc11d7bf;
    312: T0 = 32'h61b9f01f;
    313: T0 = 32'hbfc07f67;
    314: T0 = 32'h2177f80;
    315: T0 = 32'hbfbe19dc;
    316: T0 = 32'hf0006ff8;
    317: T0 = 32'h488bc09f;
    318: T0 = 32'hdf81f29f;
    319: T0 = 32'h151afe0c;
    320: T0 = 32'h7ffccf3b;
    321: T0 = 32'hf21383f8;
    322: T0 = 32'he7ff87f5;
    323: T0 = 32'hffc1ac7f;
    324: T0 = 32'h284fffff;
    325: T0 = 32'h3ffefd41;
    326: T0 = 32'he54007fe;
    327: T0 = 32'h31ffd79d;
    328: T0 = 32'hfe24c007;
    329: T0 = 32'hfedf73f3;
    330: T0 = 32'hffc7d000;
    331: T0 = 32'he81d5706;
    332: T0 = 32'he03f1409;
    333: T0 = 32'h527843ff;
    334: T0 = 32'hc90081d7;
    335: T0 = 32'hafc848ad;
    336: T0 = 32'hff009bab;
    337: T0 = 32'h3878ec9d;
    338: T0 = 32'hf66f12ff;
    339: T0 = 32'h280379fd;
    340: T0 = 32'h6db566c9;
    341: T0 = 32'h530c4e92;
    342: T0 = 32'haa0712f0;
    343: T0 = 32'hf9e8e3ea;
    344: T0 = 32'he70f80cb;
    345: T0 = 32'h14a05654;
    346: T0 = 32'h4ae916d7;
    347: T0 = 32'h1d4c380a;
    348: T0 = 32'h4bd13029;
    349: T0 = 32'h3005a40;
    350: T0 = 32'h180000fd;
    351: T0 = 32'h9f3f8;
    352: T0 = 32'h6c40fd0a;
    353: T0 = 32'h1f83f01f;
    354: T0 = 32'h8e54f805;
    355: T0 = 32'hb8ff2713;
    356: T0 = 32'hfeaf8e00;
    357: T0 = 32'hd57f01e1;
    358: T0 = 32'hdff3b0f8;
    359: T0 = 32'ha3dff10b;
    360: T0 = 32'hfeff208f;
    361: T0 = 32'hfb7f87fe;
    362: T0 = 32'hfffffcf9;
    363: T0 = 32'h9bd7303f;
    364: T0 = 32'hff7f3ff2;
    365: T0 = 32'he01d7001;
    366: T0 = 32'hffe001f7;
    367: T0 = 32'h1e6c0;
    368: T0 = 32'h1f3c7f0e;
    369: T0 = 32'hd0006ab8;
    370: T0 = 32'h641cff0;
    371: T0 = 32'h16008324;
    372: T0 = 32'h3e717c;
    373: T0 = 32'hc408d01c;
    374: T0 = 32'h8006c243;
    375: T0 = 32'h65c03d03;
    376: T0 = 32'h101580;
    377: T0 = 32'h3ca0a382;
    378: T0 = 32'h19327;
    379: T0 = 32'h4fee1a27;
    380: T0 = 32'habdedf3;
    381: T0 = 32'hfefe0721;
    382: T0 = 32'he1bf1dfe;
    383: T0 = 32'hffffc048;
    384: T0 = 32'hfd0830df;
    385: T0 = 32'hb5ff8847;
    386: T0 = 32'hf3e22801;
    387: T0 = 32'hba730001;
    388: T0 = 32'h20055922;
    389: T0 = 32'h8d330009;
    390: T0 = 32'h383aca4;
    391: T0 = 32'hb6777a99;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T5 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T6 = reset ? 1'h0 : restartRegs_0;
  assign T7 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_8(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T5;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T6;
  reg  restartRegs_0;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (addr)
    0: T0 = 32'he836ff9b;
    1: T0 = 32'h1db7d819;
    2: T0 = 32'h96787a21;
    3: T0 = 32'ha98a4a78;
    4: T0 = 32'h2d5c2ff5;
    5: T0 = 32'hb72a9f94;
    6: T0 = 32'hf7a0187f;
    7: T0 = 32'hb201fe13;
    8: T0 = 32'h1e22e405;
    9: T0 = 32'hb0fcfffe;
    10: T0 = 32'he7afd121;
    11: T0 = 32'hcf4f3ffc;
    12: T0 = 32'hfe3f0572;
    13: T0 = 32'hfa977fff;
    14: T0 = 32'h97e08028;
    15: T0 = 32'h1229ffff;
    16: T0 = 32'h677ff800;
    17: T0 = 32'hf0c1023f;
    18: T0 = 32'h28fdff00;
    19: T0 = 32'h2f8700f3;
    20: T0 = 32'h805b8c80;
    21: T0 = 32'hf038000a;
    22: T0 = 32'h7a02dd10;
    23: T0 = 32'hdf010188;
    24: T0 = 32'h13c4ac48;
    25: T0 = 32'ha9f8001f;
    26: T0 = 32'h80f87740;
    27: T0 = 32'h837d8a00;
    28: T0 = 32'hdb8307f4;
    29: T0 = 32'h3e2fec00;
    30: T0 = 32'hc5dc300f;
    31: T0 = 32'he1f7f840;
    32: T0 = 32'hec5f0b83;
    33: T0 = 32'hea1fffa4;
    34: T0 = 32'hfdaf007f;
    35: T0 = 32'hf10bfbc;
    36: T0 = 32'hff1fa57;
    37: T0 = 32'h4f5fce3;
    38: T0 = 32'h40ffd89e;
    39: T0 = 32'hebcfffe5;
    40: T0 = 32'h7f0fbf9d;
    41: T0 = 32'hfe1fcfff;
    42: T0 = 32'hd71f706c;
    43: T0 = 32'h17e2727e;
    44: T0 = 32'h7fc00001;
    45: T0 = 32'h20cf8fe;
    46: T0 = 32'h96f06e01;
    47: T0 = 32'hc846599f;
    48: T0 = 32'hc134f641;
    49: T0 = 32'h4439d4f4;
    50: T0 = 32'hb4c66bb0;
    51: T0 = 32'h123171d9;
    52: T0 = 32'h6bc2d8c5;
    53: T0 = 32'h11b82992;
    54: T0 = 32'he6fd0ae2;
    55: T0 = 32'h1c8a1600;
    56: T0 = 32'h30001021;
    57: T0 = 32'h49d7f22;
    58: T0 = 32'h6d00fc05;
    59: T0 = 32'hfffe43eb;
    60: T0 = 32'h81f6ff00;
    61: T0 = 32'he9ff19e9;
    62: T0 = 32'h476cb440;
    63: T0 = 32'hfc010466;
    64: T0 = 32'he861800;
    65: T0 = 32'h47d000d1;
    66: T0 = 32'h8030a380;
    67: T0 = 32'h2b7e001b;
    68: T0 = 32'hfb12fb54;
    69: T0 = 32'hfedf0001;
    70: T0 = 32'h7c8f1d4c;
    71: T0 = 32'hfff04200;
    72: T0 = 32'h6ba9c1fc;
    73: T0 = 32'hbffec438;
    74: T0 = 32'he3aabf1e;
    75: T0 = 32'h3f1fa27;
    76: T0 = 32'hc0b037f9;
    77: T0 = 32'h5fcea1;
    78: T0 = 32'hf8078fff;
    79: T0 = 32'h7b01fc65;
    80: T0 = 32'h700f07f;
    81: T0 = 32'ha90ffc7;
    82: T0 = 32'h80003f23;
    83: T0 = 32'h202ffc;
    84: T0 = 32'hb8000db4;
    85: T0 = 32'h1eddf8b;
    86: T0 = 32'he56000df;
    87: T0 = 32'h4cffd4ba;
    88: T0 = 32'hed070000;
    89: T0 = 32'h7fff8b2d;
    90: T0 = 32'hf5b11001;
    91: T0 = 32'hb5ff01e8;
    92: T0 = 32'hf40fad00;
    93: T0 = 32'hbebf0000;
    94: T0 = 32'h900051a8;
    95: T0 = 32'hb3e501a;
    96: T0 = 32'h8400ce2e;
    97: T0 = 32'hc3ccd0cf;
    98: T0 = 32'hd71a93e5;
    99: T0 = 32'h90b2fe1e;
    100: T0 = 32'h28b1517b;
    101: T0 = 32'h2b18e9dd;
    102: T0 = 32'h6712f6e8;
    103: T0 = 32'h41a50d42;
    104: T0 = 32'h65058180;
    105: T0 = 32'hea01f8d6;
    106: T0 = 32'h7fe430dc;
    107: T0 = 32'h2f807dff;
    108: T0 = 32'hfffca0f;
    109: T0 = 32'hfd70f827;
    110: T0 = 32'h1be1dfa;
    111: T0 = 32'hefa0ed00;
    112: T0 = 32'h383e0000;
    113: T0 = 32'hf7fc0590;
    114: T0 = 32'ha9030000;
    115: T0 = 32'h3f0f079d;
    116: T0 = 32'h1cd07f80;
    117: T0 = 32'h3e0009b;
    118: T0 = 32'had858;
    119: T0 = 32'hb81ef80e;
    120: T0 = 32'hf002bf68;
    121: T0 = 32'h3fc08ff9;
    122: T0 = 32'h1e00f4f9;
    123: T0 = 32'hffffeff;
    124: T0 = 32'hf8cc7fd3;
    125: T0 = 32'hb0d75bdf;
    126: T0 = 32'hbfcef3fd;
    127: T0 = 32'h7f8564ff;
    128: T0 = 32'h86ff3f0f;
    129: T0 = 32'he63e7ee0;
    130: T0 = 32'hc46f0020;
    131: T0 = 32'hfa22029e;
    132: T0 = 32'h413a000;
    133: T0 = 32'h6f000016;
    134: T0 = 32'h223fc00;
    135: T0 = 32'h3803006;
    136: T0 = 32'hd8082fa;
    137: T0 = 32'h5e0ff80;
    138: T0 = 32'h1ce7a57;
    139: T0 = 32'he0d3b7ff;
    140: T0 = 32'hc013fc1a;
    141: T0 = 32'h1205938a;
    142: T0 = 32'hf8230004;
    143: T0 = 32'h4fda2c50;
    144: T0 = 32'hed941000;
    145: T0 = 32'ha5917547;
    146: T0 = 32'h1ea1d52b;
    147: T0 = 32'h7940007f;
    148: T0 = 32'h4bbf6370;
    149: T0 = 32'ha86591a4;
    150: T0 = 32'h1c01f5fe;
    151: T0 = 32'hdcf57242;
    152: T0 = 32'h36dc05d4;
    153: T0 = 32'h3b29c00;
    154: T0 = 32'h2f000019;
    155: T0 = 32'h30e5c0;
    156: T0 = 32'h92f40407;
    157: T0 = 32'ha003ee60;
    158: T0 = 32'h31af07c0;
    159: T0 = 32'hf800023c;
    160: T0 = 32'h373c0fc;
    161: T0 = 32'hfff0e366;
    162: T0 = 32'h38349c07;
    163: T0 = 32'hc7eb7c7f;
    164: T0 = 32'h3c1e8d0;
    165: T0 = 32'h57e23cf;
    166: T0 = 32'hc07cff28;
    167: T0 = 32'he0f7c738;
    168: T0 = 32'h380f0ff9;
    169: T0 = 32'hfe07e3bf;
    170: T0 = 32'ha401f87f;
    171: T0 = 32'h3fe0f94f;
    172: T0 = 32'hda05f81;
    173: T0 = 32'h3fc0190;
    174: T0 = 32'h1c0407a;
    175: T0 = 32'h401ef02b;
    176: T0 = 32'he8309a07;
    177: T0 = 32'h50000f00;
    178: T0 = 32'h6e20fa0;
    179: T0 = 32'hd5400078;
    180: T0 = 32'h65e8126;
    181: T0 = 32'ha032c007;
    182: T0 = 32'h80977802;
    183: T0 = 32'h89043c00;
    184: T0 = 32'h900869c0;
    185: T0 = 32'h21800fe0;
    186: T0 = 32'h8c095e0;
    187: T0 = 32'h33b19c7;
    188: T0 = 32'hc0461ffe;
    189: T0 = 32'hd0378171;
    190: T0 = 32'hc080ea7f;
    191: T0 = 32'h57c1680c;
    192: T0 = 32'h1585e3ab;
    193: T0 = 32'hd370ffee;
    194: T0 = 32'h15cc735a;
    195: T0 = 32'hcae2a89e;
    196: T0 = 32'hb56a84a6;
    197: T0 = 32'h7b824c5c;
    198: T0 = 32'h3bb45270;
    199: T0 = 32'h98d793c1;
    200: T0 = 32'hba8ecc3d;
    201: T0 = 32'h27ffa8ff;
    202: T0 = 32'hce1e66c1;
    203: T0 = 32'h9abf1ef8;
    204: T0 = 32'hff8c232e;
    205: T0 = 32'h240ff0fe;
    206: T0 = 32'hffe2dcc2;
    207: T0 = 32'h5863f83;
    208: T0 = 32'hdf0039ad;
    209: T0 = 32'hcc3f8;
    210: T0 = 32'hdfc087c6;
    211: T0 = 32'h83c0f;
    212: T0 = 32'h61fc787e;
    213: T0 = 32'he00bef40;
    214: T0 = 32'h10fd0387;
    215: T0 = 32'he00034b3;
    216: T0 = 32'hfa9e8b3c;
    217: T0 = 32'h4407e015;
    218: T0 = 32'h7ffae8f3;
    219: T0 = 32'hf9e0ff00;
    220: T0 = 32'h9ff023f;
    221: T0 = 32'hfe4ffff8;
    222: T0 = 32'h702fe166;
    223: T0 = 32'h1fa0c0ff;
    224: T0 = 32'h963f40;
    225: T0 = 32'h647a3803;
    226: T0 = 32'h5a0413fc;
    227: T0 = 32'h41fc7f40;
    228: T0 = 32'h80c0833f;
    229: T0 = 32'h97ffd15;
    230: T0 = 32'hfc64d9a1;
    231: T0 = 32'h207f9ec8;
    232: T0 = 32'hffc56ec0;
    233: T0 = 32'h34ff000f;
    234: T0 = 32'hfe1e87fc;
    235: T0 = 32'hc68fe010;
    236: T0 = 32'h7fff9704;
    237: T0 = 32'he03a0f41;
    238: T0 = 32'hcfff341c;
    239: T0 = 32'hc00219fd;
    240: T0 = 32'h3c7f3f01;
    241: T0 = 32'hfc805cf9;
    242: T0 = 32'h1bf6c04b;
    243: T0 = 32'h5029de09;
    244: T0 = 32'h43908ddd;
    245: T0 = 32'hf80df1c9;
    246: T0 = 32'hed83e0d3;
    247: T0 = 32'he8d7d1a4;
    248: T0 = 32'hf2d1b19e;
    249: T0 = 32'h9a238002;
    250: T0 = 32'h585302b3;
    251: T0 = 32'h949a5f60;
    252: T0 = 32'hdbc0fa1a;
    253: T0 = 32'h7d5a47f;
    254: T0 = 32'he9e0ffe9;
    255: T0 = 32'h807f19b7;
    256: T0 = 32'hc87efffe;
    257: T0 = 32'h907b00a7;
    258: T0 = 32'hbfd3fffe;
    259: T0 = 32'heb87def2;
    260: T0 = 32'h1ff887ff;
    261: T0 = 32'hcf001c0f;
    262: T0 = 32'h381e74ff;
    263: T0 = 32'h30f68069;
    264: T0 = 32'h8383018b;
    265: T0 = 32'hec7f4007;
    266: T0 = 32'h207d720c;
    267: T0 = 32'hdf9b2c20;
    268: T0 = 32'h28070737;
    269: T0 = 32'h13ebcd00;
    270: T0 = 32'h2000070;
    271: T0 = 32'hb81d008;
    272: T0 = 32'h4f00007;
    273: T0 = 32'h2be3000;
    274: T0 = 32'h601da000;
    275: T0 = 32'h18020143;
    276: T0 = 32'h37037b64;
    277: T0 = 32'h3d00fc00;
    278: T0 = 32'h1b787fc9;
    279: T0 = 32'h80e0dff1;
    280: T0 = 32'h177fffd;
    281: T0 = 32'hf81de5ff;
    282: T0 = 32'h600fffff;
    283: T0 = 32'hff89ee7f;
    284: T0 = 32'h168ffff;
    285: T0 = 32'hffe1f89a;
    286: T0 = 32'h1f822fff;
    287: T0 = 32'hf7fcf810;
    288: T0 = 32'hc0f36187;
    289: T0 = 32'h5bff7210;
    290: T0 = 32'hfe6d8260;
    291: T0 = 32'h23974a81;
    292: T0 = 32'h1ba29671;
    293: T0 = 32'h71149502;
    294: T0 = 32'h88018fbd;
    295: T0 = 32'h4eeeb00;
    296: T0 = 32'h23de2e6e;
    297: T0 = 32'h2ec14907;
    298: T0 = 32'h27b807e7;
    299: T0 = 32'h2174dbbc;
    300: T0 = 32'hb854e838;
    301: T0 = 32'h3fdfa6;
    302: T0 = 32'hff8f5207;
    303: T0 = 32'h781b7fff;
    304: T0 = 32'h1cbfe1a2;
    305: T0 = 32'h76c009f7;
    306: T0 = 32'h3fdf94;
    307: T0 = 32'hfdc88402;
    308: T0 = 32'h4071efb;
    309: T0 = 32'hdfdf1908;
    310: T0 = 32'h18cf01e3;
    311: T0 = 32'hfedef008;
    312: T0 = 32'hfb77e00f;
    313: T0 = 32'hffe0f479;
    314: T0 = 32'hf8bbe00;
    315: T0 = 32'h3ffc0ff0;
    316: T0 = 32'h7d0bfe;
    317: T0 = 32'hcff8f0ff;
    318: T0 = 32'h7e31f;
    319: T0 = 32'h7d7ff3ff;
    320: T0 = 32'hfc00fbb3;
    321: T0 = 32'h79bde13;
    322: T0 = 32'hbf84bfe8;
    323: T0 = 32'h20f829e1;
    324: T0 = 32'heff013ff;
    325: T0 = 32'he1fe85f;
    326: T0 = 32'hd47ff03f;
    327: T0 = 32'hf027ff6b;
    328: T0 = 32'h7e975f8b;
    329: T0 = 32'hf861e7d;
    330: T0 = 32'h1f8ef9fd;
    331: T0 = 32'h80f8e0ce;
    332: T0 = 32'hf8fe493f;
    333: T0 = 32'h407fff31;
    334: T0 = 32'hfb020058;
    335: T0 = 32'h281ff3;
    336: T0 = 32'hb700d80b;
    337: T0 = 32'h400d56ff;
    338: T0 = 32'hb1f86005;
    339: T0 = 32'h7ff0d85e;
    340: T0 = 32'hbf56a877;
    341: T0 = 32'hbb7f9adb;
    342: T0 = 32'h313183d2;
    343: T0 = 32'hb17a2f60;
    344: T0 = 32'h5fc84e14;
    345: T0 = 32'hfc61019e;
    346: T0 = 32'ha70c8b1e;
    347: T0 = 32'hc1f8f043;
    348: T0 = 32'h278f0a78;
    349: T0 = 32'hbf92b480;
    350: T0 = 32'hdfc101ad;
    351: T0 = 32'hf7bf6f0;
    352: T0 = 32'hb3ecf580;
    353: T0 = 32'h83df34fe;
    354: T0 = 32'hf07edf00;
    355: T0 = 32'hc03b52b5;
    356: T0 = 32'hf1775f0;
    357: T0 = 32'h380705fd;
    358: T0 = 32'h7ffbcecf;
    359: T0 = 32'habc0f83c;
    360: T0 = 32'h7ff4605;
    361: T0 = 32'hfc30bfc2;
    362: T0 = 32'h7f01cd;
    363: T0 = 32'hef8ea2fe;
    364: T0 = 32'he007f004;
    365: T0 = 32'hfb3af60d;
    366: T0 = 32'hde0f8780;
    367: T0 = 32'h7f8816c0;
    368: T0 = 32'h1d6107fc;
    369: T0 = 32'h937ac1ee;
    370: T0 = 32'ha06e387f;
    371: T0 = 32'h38bff80a;
    372: T0 = 32'hfa08e7c3;
    373: T0 = 32'hd7f91fa0;
    374: T0 = 32'h7f9dfaf0;
    375: T0 = 32'hc05d40ff;
    376: T0 = 32'ha7cbeff3;
    377: T0 = 32'h93bf603;
    378: T0 = 32'hf8bc3fdb;
    379: T0 = 32'hc2b041f8;
    380: T0 = 32'h3f2fc1cd;
    381: T0 = 32'hfc75b49e;
    382: T0 = 32'h35db01e;
    383: T0 = 32'h7f84fee9;
    384: T0 = 32'h20356250;
    385: T0 = 32'hbff803f7;
    386: T0 = 32'h831dcc80;
    387: T0 = 32'h25df0878;
    388: T0 = 32'hfc01d138;
    389: T0 = 32'h4975c146;
    390: T0 = 32'h8fc1f6bd;
    391: T0 = 32'hb626b3df;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T5 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T6 = reset ? 1'h0 : restartRegs_0;
  assign T7 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_9(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T5;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T6;
  reg  restartRegs_0;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (addr)
    0: T0 = 32'heb2eab67;
    1: T0 = 32'hcdfbfd75;
    2: T0 = 32'ha03a72ee;
    3: T0 = 32'h37c68185;
    4: T0 = 32'hfd004224;
    5: T0 = 32'hde3e02e9;
    6: T0 = 32'hbe27731e;
    7: T0 = 32'h4fffe071;
    8: T0 = 32'hfff33078;
    9: T0 = 32'h50ff0f81;
    10: T0 = 32'hf8f40e4f;
    11: T0 = 32'hcec3e870;
    12: T0 = 32'h11efc129;
    13: T0 = 32'hff8837cf;
    14: T0 = 32'h5790f;
    15: T0 = 32'h3e78db14;
    16: T0 = 32'h48000398;
    17: T0 = 32'h4078800;
    18: T0 = 32'h3c40003f;
    19: T0 = 32'he0feb8;
    20: T0 = 32'heee001;
    21: T0 = 32'h911e0ff6;
    22: T0 = 32'he01e840e;
    23: T0 = 32'hff97f0ff;
    24: T0 = 32'h5e00fc01;
    25: T0 = 32'h173e3f0d;
    26: T0 = 32'hfde06efc;
    27: T0 = 32'h3941f0;
    28: T0 = 32'h9fff82ba;
    29: T0 = 32'hf8092617;
    30: T0 = 32'haf7e7c23;
    31: T0 = 32'he780f701;
    32: T0 = 32'h4aff09c0;
    33: T0 = 32'hbe4e0f63;
    34: T0 = 32'hf383709c;
    35: T0 = 32'h7d0ae07f;
    36: T0 = 32'h5ffb7d0b;
    37: T0 = 32'haaa15e17;
    38: T0 = 32'h3fff71f3;
    39: T0 = 32'hffb59fe8;
    40: T0 = 32'h1e06419a;
    41: T0 = 32'h6f3db1fe;
    42: T0 = 32'h40000035;
    43: T0 = 32'h5ff34adf;
    44: T0 = 32'h39017c25;
    45: T0 = 32'h17801a4f;
    46: T0 = 32'hd625d1f5;
    47: T0 = 32'h988a6386;
    48: T0 = 32'hd455c1e0;
    49: T0 = 32'hb856dfc7;
    50: T0 = 32'hfffe427a;
    51: T0 = 32'h964c39f8;
    52: T0 = 32'h74df6ce8;
    53: T0 = 32'hf5fbe9a2;
    54: T0 = 32'h240da325;
    55: T0 = 32'hbc43dffe;
    56: T0 = 32'h2000e01b;
    57: T0 = 32'hbeb5c2ec;
    58: T0 = 32'h3a00f758;
    59: T0 = 32'hffd700bf;
    60: T0 = 32'h7de8ff07;
    61: T0 = 32'hffe8ca2f;
    62: T0 = 32'heafc7ff;
    63: T0 = 32'hf780fde9;
    64: T0 = 32'hf8000a;
    65: T0 = 32'h2fff0f02;
    66: T0 = 32'he8bf2fc0;
    67: T0 = 32'hf9ff0000;
    68: T0 = 32'hf2ff0000;
    69: T0 = 32'h7eef0000;
    70: T0 = 32'hff0e0007;
    71: T0 = 32'h61fa2600;
    72: T0 = 32'hb7e00400;
    73: T0 = 32'h60308f0;
    74: T0 = 32'h3afe01e1;
    75: T0 = 32'he0601c56;
    76: T0 = 32'h79f723e;
    77: T0 = 32'h7e07ee70;
    78: T0 = 32'h707d7f63;
    79: T0 = 32'h87f01fef;
    80: T0 = 32'h830f16fc;
    81: T0 = 32'hf85f91f7;
    82: T0 = 32'hfc23f8a3;
    83: T0 = 32'h7e4f5f0f;
    84: T0 = 32'h3ffef39d;
    85: T0 = 32'haff509e8;
    86: T0 = 32'hfeff87f3;
    87: T0 = 32'hfcfee57c;
    88: T0 = 32'hdfd3de1f;
    89: T0 = 32'h5ffb7e0d;
    90: T0 = 32'hc350cf80;
    91: T0 = 32'hf1ff0224;
    92: T0 = 32'hfe000720;
    93: T0 = 32'h918f0007;
    94: T0 = 32'h6100bd38;
    95: T0 = 32'h32c89011;
    96: T0 = 32'ha05929bb;
    97: T0 = 32'h7741688e;
    98: T0 = 32'h1e078b7b;
    99: T0 = 32'h489e4755;
    100: T0 = 32'hc2765222;
    101: T0 = 32'hdbb5a77d;
    102: T0 = 32'h5244407d;
    103: T0 = 32'hfbd8ff0f;
    104: T0 = 32'h1108946f;
    105: T0 = 32'hdffeffe3;
    106: T0 = 32'hc8249cff;
    107: T0 = 32'h2362fe03;
    108: T0 = 32'h3d024dff;
    109: T0 = 32'h103dd040;
    110: T0 = 32'hffd00534;
    111: T0 = 32'he0470000;
    112: T0 = 32'hffff0025;
    113: T0 = 32'hffcf5a00;
    114: T0 = 32'h13ff0188;
    115: T0 = 32'hffb42a0;
    116: T0 = 32'h15b00061;
    117: T0 = 32'h7f0347;
    118: T0 = 32'h400e8e;
    119: T0 = 32'h8000c01a;
    120: T0 = 32'h4ed36;
    121: T0 = 32'h1300ae00;
    122: T0 = 32'h60000a10;
    123: T0 = 32'h1e4014e0;
    124: T0 = 32'h1fc400fa;
    125: T0 = 32'h168b64f;
    126: T0 = 32'h11fcec51;
    127: T0 = 32'hc00d3fe9;
    128: T0 = 32'h390edcff;
    129: T0 = 32'hcc00fe39;
    130: T0 = 32'h9c41ffff;
    131: T0 = 32'h1de0ff9f;
    132: T0 = 32'h7acbeff;
    133: T0 = 32'ha1defffd;
    134: T0 = 32'hf0fbafab;
    135: T0 = 32'h907dfffc;
    136: T0 = 32'h7f400f7f;
    137: T0 = 32'h2cfce0e;
    138: T0 = 32'hfacc0149;
    139: T0 = 32'h8090e200;
    140: T0 = 32'h4fdb0035;
    141: T0 = 32'h38bec70;
    142: T0 = 32'hcabc0005;
    143: T0 = 32'h6bb8d80d;
    144: T0 = 32'hb5b4c41;
    145: T0 = 32'he28b9586;
    146: T0 = 32'had372eb3;
    147: T0 = 32'h4042710f;
    148: T0 = 32'hb28a29cc;
    149: T0 = 32'h5ead654d;
    150: T0 = 32'h10a6a6a2;
    151: T0 = 32'hf3db17c8;
    152: T0 = 32'hfe960047;
    153: T0 = 32'heb2cc800;
    154: T0 = 32'h47ffc851;
    155: T0 = 32'h27b880e6;
    156: T0 = 32'h65fffb00;
    157: T0 = 32'hc00f1567;
    158: T0 = 32'haedfffc2;
    159: T0 = 32'hc80f874;
    160: T0 = 32'h3523fff;
    161: T0 = 32'h401cffc0;
    162: T0 = 32'he65ff;
    163: T0 = 32'hed00e3fe;
    164: T0 = 32'hfd3f;
    165: T0 = 32'hfffe3f;
    166: T0 = 32'hfc00ff88;
    167: T0 = 32'h1fba6e0;
    168: T0 = 32'hffe807c1;
    169: T0 = 32'hf7fd24de;
    170: T0 = 32'he8bfc000;
    171: T0 = 32'h7fff2111;
    172: T0 = 32'hfe800200;
    173: T0 = 32'h1fff0b9;
    174: T0 = 32'hffe4803b;
    175: T0 = 32'h400fffc3;
    176: T0 = 32'hfff81403;
    177: T0 = 32'he4007ffe;
    178: T0 = 32'hfff4280;
    179: T0 = 32'h9b001087;
    180: T0 = 32'h19ff0ce8;
    181: T0 = 32'h83a2f9c0;
    182: T0 = 32'hc0fc0004;
    183: T0 = 32'hc00ba3eb;
    184: T0 = 32'ha23f8000;
    185: T0 = 32'hfd811c1f;
    186: T0 = 32'h24c9fff9;
    187: T0 = 32'h5d00892b;
    188: T0 = 32'hd237ff;
    189: T0 = 32'hb7c0fffb;
    190: T0 = 32'h6345bd3;
    191: T0 = 32'h91ffbfff;
    192: T0 = 32'hb730d296;
    193: T0 = 32'h2f570376;
    194: T0 = 32'h4818d820;
    195: T0 = 32'h48c8a97a;
    196: T0 = 32'hf982cb94;
    197: T0 = 32'h667567ef;
    198: T0 = 32'h4dbf45b1;
    199: T0 = 32'h51168a02;
    200: T0 = 32'hd429f00c;
    201: T0 = 32'h45a2ce7c;
    202: T0 = 32'hd059c200;
    203: T0 = 32'h3bf50c80;
    204: T0 = 32'hffa06680;
    205: T0 = 32'h837f804c;
    206: T0 = 32'hfbfce59c;
    207: T0 = 32'h430f683f;
    208: T0 = 32'hffdbff2d;
    209: T0 = 32'h107c4ae7;
    210: T0 = 32'h80beffaf;
    211: T0 = 32'hbb75555b;
    212: T0 = 32'h60001ffd;
    213: T0 = 32'hd00148;
    214: T0 = 32'h8e830060;
    215: T0 = 32'h1e0f0008;
    216: T0 = 32'h98740000;
    217: T0 = 32'h1ff0001;
    218: T0 = 32'hff020580;
    219: T0 = 32'h50070000;
    220: T0 = 32'h7fd00178;
    221: T0 = 32'h10e003;
    222: T0 = 32'h3f84cf7;
    223: T0 = 32'h80cfbf04;
    224: T0 = 32'hbc0745e7;
    225: T0 = 32'h300f3bf8;
    226: T0 = 32'hfb748000;
    227: T0 = 32'hf00104ff;
    228: T0 = 32'h77437c00;
    229: T0 = 32'h3b80001a;
    230: T0 = 32'h79a0500;
    231: T0 = 32'h6378c000;
    232: T0 = 32'h1f35843;
    233: T0 = 32'h80147fc2;
    234: T0 = 32'hc271f601;
    235: T0 = 32'h44f1cfff;
    236: T0 = 32'h178ff1a;
    237: T0 = 32'hff6ea93f;
    238: T0 = 32'he07f7ff8;
    239: T0 = 32'hffb4b942;
    240: T0 = 32'h6c0749bf;
    241: T0 = 32'h37fee9a6;
    242: T0 = 32'had40876f;
    243: T0 = 32'hd6ff7883;
    244: T0 = 32'hf9484fc0;
    245: T0 = 32'hdc6f3be7;
    246: T0 = 32'hc49d08f;
    247: T0 = 32'h71c55ca8;
    248: T0 = 32'hccb39dc4;
    249: T0 = 32'h4636fea3;
    250: T0 = 32'h48cb25b6;
    251: T0 = 32'h6c1a62f0;
    252: T0 = 32'hd4c30172;
    253: T0 = 32'h3fa50e78;
    254: T0 = 32'h44ff000b;
    255: T0 = 32'ha7fc18ce;
    256: T0 = 32'ha85f0000;
    257: T0 = 32'h1a770064;
    258: T0 = 32'hfe29800e;
    259: T0 = 32'h9ff70003;
    260: T0 = 32'hff3b6400;
    261: T0 = 32'h7df0000;
    262: T0 = 32'hff06a770;
    263: T0 = 32'hbf8083;
    264: T0 = 32'h3f77;
    265: T0 = 32'h1afefc;
    266: T0 = 32'hb000f7fd;
    267: T0 = 32'h415e7ef;
    268: T0 = 32'hc809fff;
    269: T0 = 32'h60edff;
    270: T0 = 32'hf500ffff;
    271: T0 = 32'h3fe91;
    272: T0 = 32'h3fc41ff7;
    273: T0 = 32'hc100fff2;
    274: T0 = 32'h3f1b577;
    275: T0 = 32'h90008fff;
    276: T0 = 32'h8000e2c0;
    277: T0 = 32'h16104ff;
    278: T0 = 32'hd000e8f0;
    279: T0 = 32'h6c003;
    280: T0 = 32'hcf700800;
    281: T0 = 32'hf0005c02;
    282: T0 = 32'hfc7f1801;
    283: T0 = 32'hfffe1bf0;
    284: T0 = 32'hfbaf0000;
    285: T0 = 32'hffff03b6;
    286: T0 = 32'hff162000;
    287: T0 = 32'h4ff7000e;
    288: T0 = 32'h2ff0eff6;
    289: T0 = 32'hac10a2f7;
    290: T0 = 32'hffff1a67;
    291: T0 = 32'ha9e7704a;
    292: T0 = 32'hfdb1b02;
    293: T0 = 32'h8e90e39a;
    294: T0 = 32'h3a9c2eb7;
    295: T0 = 32'hdcb4de5;
    296: T0 = 32'hb9e86d67;
    297: T0 = 32'hb149412f;
    298: T0 = 32'h4540f643;
    299: T0 = 32'h7fbd1fad;
    300: T0 = 32'h728ebe78;
    301: T0 = 32'h440c465;
    302: T0 = 32'h5b7b1ff;
    303: T0 = 32'hfb43f8ff;
    304: T0 = 32'h59cc23;
    305: T0 = 32'h85001f21;
    306: T0 = 32'h470bfe44;
    307: T0 = 32'hbc44807d;
    308: T0 = 32'h42b79db8;
    309: T0 = 32'h8ab85403;
    310: T0 = 32'h3406385e;
    311: T0 = 32'h387d4748;
    312: T0 = 32'h79e1c7eb;
    313: T0 = 32'hf80ff44;
    314: T0 = 32'h2817fff;
    315: T0 = 32'h953cbffd;
    316: T0 = 32'he00291ff;
    317: T0 = 32'h5007f87e;
    318: T0 = 32'hfff8eadf;
    319: T0 = 32'h8838fd01;
    320: T0 = 32'h9fff10fc;
    321: T0 = 32'hf060af08;
    322: T0 = 32'ha0ff0c86;
    323: T0 = 32'hfc047c60;
    324: T0 = 32'hb80701e8;
    325: T0 = 32'h18008208;
    326: T0 = 32'h1480403e;
    327: T0 = 32'he324;
    328: T0 = 32'h1ec0003;
    329: T0 = 32'ha0087c89;
    330: T0 = 32'h380200;
    331: T0 = 32'hc8081fec;
    332: T0 = 32'h206fc340;
    333: T0 = 32'hff20bfff;
    334: T0 = 32'h800ff844;
    335: T0 = 32'h3fc2cffb;
    336: T0 = 32'hb003c00d;
    337: T0 = 32'h4ff137e;
    338: T0 = 32'h9400fe17;
    339: T0 = 32'h27360159;
    340: T0 = 32'h9d8015ff;
    341: T0 = 32'hac5e141c;
    342: T0 = 32'hac05a6cc;
    343: T0 = 32'hb5bf2882;
    344: T0 = 32'hf2fa93c6;
    345: T0 = 32'h3b556258;
    346: T0 = 32'h79a72f22;
    347: T0 = 32'ha4ec7a32;
    348: T0 = 32'h20a0ff02;
    349: T0 = 32'h3bcf13f;
    350: T0 = 32'h10fcbec6;
    351: T0 = 32'h804f4f49;
    352: T0 = 32'ha4befffc;
    353: T0 = 32'ha800fc1f;
    354: T0 = 32'hce65ffff;
    355: T0 = 32'hc005ffb7;
    356: T0 = 32'h2824beff;
    357: T0 = 32'h1c00000c;
    358: T0 = 32'ha5e501;
    359: T0 = 32'hfbf80001;
    360: T0 = 32'hfff13a00;
    361: T0 = 32'hd2d70000;
    362: T0 = 32'hffff01a4;
    363: T0 = 32'hfeb190f0;
    364: T0 = 32'hafff8038;
    365: T0 = 32'hff80843f;
    366: T0 = 32'h5649f280;
    367: T0 = 32'hffff1f83;
    368: T0 = 32'hc8310690;
    369: T0 = 32'h9ffe01a4;
    370: T0 = 32'hfcbfe0f2;
    371: T0 = 32'h3cff801f;
    372: T0 = 32'hffdecc10;
    373: T0 = 32'h8fd74803;
    374: T0 = 32'h7ffffb00;
    375: T0 = 32'hfd1fffc0;
    376: T0 = 32'h4bffffc7;
    377: T0 = 32'hff7697bf;
    378: T0 = 32'h90877ff8;
    379: T0 = 32'hf1a99f7;
    380: T0 = 32'h7900f3ff;
    381: T0 = 32'h1ffff;
    382: T0 = 32'h5a0ff43;
    383: T0 = 32'h5000b6ce;
    384: T0 = 32'h881fed;
    385: T0 = 32'h783fd60c;
    386: T0 = 32'h9042ff3;
    387: T0 = 32'ha7b8fc00;
    388: T0 = 32'ha570;
    389: T0 = 32'he4104386;
    390: T0 = 32'h483e5953;
    391: T0 = 32'he81ae834;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T5 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T6 = reset ? 1'h0 : restartRegs_0;
  assign T7 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_10(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T5;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T6;
  reg  restartRegs_0;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (addr)
    0: T0 = 32'h89715a2;
    1: T0 = 32'h73c94b8b;
    2: T0 = 32'h46dabfab;
    3: T0 = 32'h27e529a1;
    4: T0 = 32'hedb0bb41;
    5: T0 = 32'hb407001d;
    6: T0 = 32'hfe7c2800;
    7: T0 = 32'h1fc0005e;
    8: T0 = 32'h3fe4dc00;
    9: T0 = 32'h9af03fae;
    10: T0 = 32'h3fe0d06;
    11: T0 = 32'hd93e0028;
    12: T0 = 32'hc0fb8408;
    13: T0 = 32'h80cfd000;
    14: T0 = 32'hfe0f017c;
    15: T0 = 32'hf00e8be0;
    16: T0 = 32'hbfe0b03f;
    17: T0 = 32'h780f43f;
    18: T0 = 32'h919ff5ff;
    19: T0 = 32'hf07fff1b;
    20: T0 = 32'hff3ff9cf;
    21: T0 = 32'h1f87ffff;
    22: T0 = 32'h3ff6a2dc;
    23: T0 = 32'ha7fcdfff;
    24: T0 = 32'he7fffdc7;
    25: T0 = 32'hea8703fb;
    26: T0 = 32'h4a3e0d6;
    27: T0 = 32'h4eb4a03f;
    28: T0 = 32'h8008f801;
    29: T0 = 32'h45e6301;
    30: T0 = 32'h36000e00;
    31: T0 = 32'hf603e2;
    32: T0 = 32'h6806000;
    33: T0 = 32'h710f0005;
    34: T0 = 32'hf04e4c00;
    35: T0 = 32'h7df70008;
    36: T0 = 32'hed63a74e;
    37: T0 = 32'had7f047f;
    38: T0 = 32'h99a2fe16;
    39: T0 = 32'hfd8ebf;
    40: T0 = 32'hfc32fbf5;
    41: T0 = 32'h90f0d03f;
    42: T0 = 32'hbf3d05f7;
    43: T0 = 32'h1e0e06b8;
    44: T0 = 32'h6b7c245e;
    45: T0 = 32'hfff4f480;
    46: T0 = 32'h8b351aff;
    47: T0 = 32'h6dafa266;
    48: T0 = 32'h42fd3688;
    49: T0 = 32'h4e463a71;
    50: T0 = 32'hfe6b7450;
    51: T0 = 32'h1c1c4f29;
    52: T0 = 32'h63256bf5;
    53: T0 = 32'h2f126e78;
    54: T0 = 32'hda16e185;
    55: T0 = 32'hfb6b081f;
    56: T0 = 32'h280779ad;
    57: T0 = 32'hfff6de1a;
    58: T0 = 32'hc38fe3f3;
    59: T0 = 32'hbff9f76f;
    60: T0 = 32'h31a4d7e;
    61: T0 = 32'h8000cc42;
    62: T0 = 32'h577087;
    63: T0 = 32'h90001e06;
    64: T0 = 32'h137610;
    65: T0 = 32'hb90001f4;
    66: T0 = 32'ha3b0;
    67: T0 = 32'h2fe0000f;
    68: T0 = 32'h80c4feb8;
    69: T0 = 32'h7332f70;
    70: T0 = 32'hff3e07f6;
    71: T0 = 32'he021c6fd;
    72: T0 = 32'hd712e07f;
    73: T0 = 32'h5f01f99e;
    74: T0 = 32'h373de03;
    75: T0 = 32'hc7f03f89;
    76: T0 = 32'h1ef8780;
    77: T0 = 32'hf37f0bf7;
    78: T0 = 32'he0189954;
    79: T0 = 32'h7efe0c4;
    80: T0 = 32'hf0410286;
    81: T0 = 32'hcfff1e0b;
    82: T0 = 32'hff3f6199;
    83: T0 = 32'hfdeb81f0;
    84: T0 = 32'h7fff811d;
    85: T0 = 32'h7feb9f53;
    86: T0 = 32'h8bfe7802;
    87: T0 = 32'h7ffc3c3d;
    88: T0 = 32'hbfd827c0;
    89: T0 = 32'h80878dce;
    90: T0 = 32'h3f294bc;
    91: T0 = 32'h1800f077;
    92: T0 = 32'he63ff;
    93: T0 = 32'h1e30fc04;
    94: T0 = 32'h1a8ff;
    95: T0 = 32'h6c537743;
    96: T0 = 32'h601b4ed;
    97: T0 = 32'h92ea7e62;
    98: T0 = 32'hb05a1155;
    99: T0 = 32'h406d0afe;
    100: T0 = 32'hc8cffe89;
    101: T0 = 32'h2b1b59;
    102: T0 = 32'h79e3bf00;
    103: T0 = 32'h60300f32;
    104: T0 = 32'h998e3ff0;
    105: T0 = 32'hb5c10072;
    106: T0 = 32'h1fc07daf;
    107: T0 = 32'hadf2f883;
    108: T0 = 32'hfdfc0af9;
    109: T0 = 32'h2bb5fc4;
    110: T0 = 32'h3e0001a6;
    111: T0 = 32'h164bffc;
    112: T0 = 32'h4200f910;
    113: T0 = 32'h207bef;
    114: T0 = 32'hbc0007e3;
    115: T0 = 32'h3cd8;
    116: T0 = 32'h200007f;
    117: T0 = 32'hbe8c;
    118: T0 = 32'h10e40003;
    119: T0 = 32'hc00073cc;
    120: T0 = 32'h5e00;
    121: T0 = 32'h4600033c;
    122: T0 = 32'h13c03381;
    123: T0 = 32'hf9601838;
    124: T0 = 32'hfbff0b8;
    125: T0 = 32'hff038163;
    126: T0 = 32'h5fff1f8d;
    127: T0 = 32'hffc1a80a;
    128: T0 = 32'h7ff11f0;
    129: T0 = 32'hfcff85c4;
    130: T0 = 32'he33f410f;
    131: T0 = 32'hffe3ff11;
    132: T0 = 32'h2e058400;
    133: T0 = 32'h7ffe0fe1;
    134: T0 = 32'hc0744c80;
    135: T0 = 32'hfdff01fe;
    136: T0 = 32'h5002bb9d;
    137: T0 = 32'h327ccdff;
    138: T0 = 32'hea3d;
    139: T0 = 32'h19aeb9f;
    140: T0 = 32'hbe73;
    141: T0 = 32'h21eb82ff;
    142: T0 = 32'hd701ffe1;
    143: T0 = 32'h1fa1c6;
    144: T0 = 32'hee4ab9fb;
    145: T0 = 32'h101b8790;
    146: T0 = 32'h231b2c86;
    147: T0 = 32'h82deb414;
    148: T0 = 32'h8360ed3;
    149: T0 = 32'h95bf9211;
    150: T0 = 32'hadc64cd3;
    151: T0 = 32'h2f7c7035;
    152: T0 = 32'h36c0fa27;
    153: T0 = 32'h5ba35c00;
    154: T0 = 32'h8bfc0525;
    155: T0 = 32'h20670ff8;
    156: T0 = 32'h60f8e81f;
    157: T0 = 32'hc00472ff;
    158: T0 = 32'h489f6700;
    159: T0 = 32'hff801f0d;
    160: T0 = 32'hffdb040;
    161: T0 = 32'h8fff03e4;
    162: T0 = 32'hf0ba8580;
    163: T0 = 32'hb41f5eff;
    164: T0 = 32'h1f03fdde;
    165: T0 = 32'hf40ffff;
    166: T0 = 32'h3f8ffbf;
    167: T0 = 32'h81707fcf;
    168: T0 = 32'h87ff03a5;
    169: T0 = 32'hf815f000;
    170: T0 = 32'h507f0003;
    171: T0 = 32'hff000a00;
    172: T0 = 32'h2d030040;
    173: T0 = 32'h76c0017c;
    174: T0 = 32'h3444006;
    175: T0 = 32'h87e4600f;
    176: T0 = 32'h401c7800;
    177: T0 = 32'hf87e0f80;
    178: T0 = 32'hec000cc0;
    179: T0 = 32'hc4605fc;
    180: T0 = 32'he80e02c;
    181: T0 = 32'h376f7ff;
    182: T0 = 32'ha2b0ff08;
    183: T0 = 32'h4340eade;
    184: T0 = 32'h1f33fff2;
    185: T0 = 32'h58dbca5a;
    186: T0 = 32'he3a31f53;
    187: T0 = 32'h2c34c4c;
    188: T0 = 32'hfe340fff;
    189: T0 = 32'hd03bee08;
    190: T0 = 32'hffe7e57f;
    191: T0 = 32'h56001b67;
    192: T0 = 32'he7f91433;
    193: T0 = 32'h89df30a3;
    194: T0 = 32'hff4333b0;
    195: T0 = 32'h76b18f52;
    196: T0 = 32'hacddf950;
    197: T0 = 32'h6dbe3ac2;
    198: T0 = 32'h7f3e04d2;
    199: T0 = 32'h75875dcb;
    200: T0 = 32'ha481cffe;
    201: T0 = 32'h3ca1132a;
    202: T0 = 32'hac61be;
    203: T0 = 32'h19fc808f;
    204: T0 = 32'ha11d401f;
    205: T0 = 32'h8c63f000;
    206: T0 = 32'h3c008401;
    207: T0 = 32'hadd83e07;
    208: T0 = 32'he1faffc0;
    209: T0 = 32'h417383e0;
    210: T0 = 32'h5f1d0ffe;
    211: T0 = 32'he40dac3e;
    212: T0 = 32'hd3c1f0db;
    213: T0 = 32'hf001b23;
    214: T0 = 32'h16bc0f80;
    215: T0 = 32'h80f800b0;
    216: T0 = 32'hc41771f8;
    217: T0 = 32'hf8078009;
    218: T0 = 32'h3fce7207;
    219: T0 = 32'h15007980;
    220: T0 = 32'h1ff1cf2;
    221: T0 = 32'he7b07bbe;
    222: T0 = 32'hc007bf35;
    223: T0 = 32'h6f30bfdf;
    224: T0 = 32'h8d40f9fd;
    225: T0 = 32'h4265ff;
    226: T0 = 32'hb5f0fe0f;
    227: T0 = 32'h20057c1f;
    228: T0 = 32'h75460f80;
    229: T0 = 32'hf8010bdf;
    230: T0 = 32'h3f0c0050;
    231: T0 = 32'h376c0f7d;
    232: T0 = 32'h7fa3b936;
    233: T0 = 32'h894f9609;
    234: T0 = 32'h6fc0e0e3;
    235: T0 = 32'h40b70a83;
    236: T0 = 32'h5ffa5f98;
    237: T0 = 32'he0484800;
    238: T0 = 32'hfdf59477;
    239: T0 = 32'hf6044e01;
    240: T0 = 32'h2e820084;
    241: T0 = 32'hf7371040;
    242: T0 = 32'hf272d000;
    243: T0 = 32'h3aff2806;
    244: T0 = 32'h9702d60;
    245: T0 = 32'h41e1031a;
    246: T0 = 32'hb3471b08;
    247: T0 = 32'h1443b53a;
    248: T0 = 32'h2a75e0d0;
    249: T0 = 32'hfb04c001;
    250: T0 = 32'ha1e726c5;
    251: T0 = 32'hb08001;
    252: T0 = 32'h2fe0060c;
    253: T0 = 32'h159fe3;
    254: T0 = 32'h1400fce0;
    255: T0 = 32'h19f;
    256: T0 = 32'hc8d0ff80;
    257: T0 = 32'h30d9;
    258: T0 = 32'h14bb1fc0;
    259: T0 = 32'h3fe00e86;
    260: T0 = 32'he016ffc2;
    261: T0 = 32'h3fbf01f8;
    262: T0 = 32'hff00c418;
    263: T0 = 32'hbff001f;
    264: T0 = 32'he03ef5c9;
    265: T0 = 32'h7cab1001;
    266: T0 = 32'h7f003dce;
    267: T0 = 32'h2dfea30;
    268: T0 = 32'h8ff801fa;
    269: T0 = 32'h80ffeedd;
    270: T0 = 32'hf8bfd83f;
    271: T0 = 32'hfe9fffb4;
    272: T0 = 32'hfed7f803;
    273: T0 = 32'h5ff1ffea;
    274: T0 = 32'h1fe13b04;
    275: T0 = 32'heffed7fe;
    276: T0 = 32'h7fef7b9;
    277: T0 = 32'ha21ce83f;
    278: T0 = 32'h3ff95b;
    279: T0 = 32'hdc3a1e29;
    280: T0 = 32'he0039f52;
    281: T0 = 32'h7d832be3;
    282: T0 = 32'hc800c1df;
    283: T0 = 32'h700f0fe;
    284: T0 = 32'h2f0fc28;
    285: T0 = 32'h1d0e6d1;
    286: T0 = 32'h8172b7;
    287: T0 = 32'ha01e100b;
    288: T0 = 32'he31ea301;
    289: T0 = 32'hdb010000;
    290: T0 = 32'h1e0c8730;
    291: T0 = 32'h94009010;
    292: T0 = 32'h35fb0359;
    293: T0 = 32'hb4238d83;
    294: T0 = 32'h9b2d22b1;
    295: T0 = 32'hc207015a;
    296: T0 = 32'h8f7aa308;
    297: T0 = 32'h72f302fa;
    298: T0 = 32'h9e710003;
    299: T0 = 32'h6a4ff956;
    300: T0 = 32'h42337781;
    301: T0 = 32'h4bc0559d;
    302: T0 = 32'hc7e40;
    303: T0 = 32'h36f801fd;
    304: T0 = 32'h8021de20;
    305: T0 = 32'h1a6f03ff;
    306: T0 = 32'hfb80fc6e;
    307: T0 = 32'h11bb47ff;
    308: T0 = 32'h3fbbffbc;
    309: T0 = 32'h3f260e01;
    310: T0 = 32'hc7f83ffa;
    311: T0 = 32'h81f0e0c0;
    312: T0 = 32'hc03f07fe;
    313: T0 = 32'hf81f0036;
    314: T0 = 32'hfe7780f0;
    315: T0 = 32'hbfc00002;
    316: T0 = 32'h3fe480e;
    317: T0 = 32'ha6fe7000;
    318: T0 = 32'hf09e01f0;
    319: T0 = 32'he57f8f00;
    320: T0 = 32'h7f19e075;
    321: T0 = 32'hcbe33878;
    322: T0 = 32'hbdf9cf04;
    323: T0 = 32'hbffc6dc3;
    324: T0 = 32'hc83f3f72;
    325: T0 = 32'h79ef6778;
    326: T0 = 32'h1c80e0fe;
    327: T0 = 32'h9dffbb;
    328: T0 = 32'hffe03c07;
    329: T0 = 32'hd0013f3d;
    330: T0 = 32'hd1f8b7e0;
    331: T0 = 32'he94010a3;
    332: T0 = 32'h363ffcce;
    333: T0 = 32'h3918d884;
    334: T0 = 32'h82b8171d;
    335: T0 = 32'h7903200;
    336: T0 = 32'he02f0029;
    337: T0 = 32'he4fd3994;
    338: T0 = 32'h90630e2b;
    339: T0 = 32'h7ff517f1;
    340: T0 = 32'hf42d007d;
    341: T0 = 32'h49ffcd6a;
    342: T0 = 32'h327ad20d;
    343: T0 = 32'h919e1ec7;
    344: T0 = 32'h1eed7fc0;
    345: T0 = 32'h8faa3777;
    346: T0 = 32'h9011f00f;
    347: T0 = 32'h8213e7f7;
    348: T0 = 32'hfa82f866;
    349: T0 = 32'h16f713ff;
    350: T0 = 32'h5fc0fffd;
    351: T0 = 32'h830b6fff;
    352: T0 = 32'h26fcfff5;
    353: T0 = 32'h1ef12b;
    354: T0 = 32'h259bffff;
    355: T0 = 32'h600ffd6;
    356: T0 = 32'hcbe63ff;
    357: T0 = 32'hbfcdfff;
    358: T0 = 32'he3152808;
    359: T0 = 32'h283f0019;
    360: T0 = 32'hfe1c0ac3;
    361: T0 = 32'hc6d72000;
    362: T0 = 32'h7df302a0;
    363: T0 = 32'h1de70f04;
    364: T0 = 32'h9fff4031;
    365: T0 = 32'hf1f939f0;
    366: T0 = 32'h22fd8e03;
    367: T0 = 32'h41f315f;
    368: T0 = 32'hf6aef8e0;
    369: T0 = 32'he0418280;
    370: T0 = 32'h1f1f1d8e;
    371: T0 = 32'h7804621b;
    372: T0 = 32'h1f0ad98;
    373: T0 = 32'h4680c009;
    374: T0 = 32'h1f0585;
    375: T0 = 32'h92ac0f3e;
    376: T0 = 32'h41c1ffc4;
    377: T0 = 32'h723522ff;
    378: T0 = 32'h940efffc;
    379: T0 = 32'h6f41447e;
    380: T0 = 32'h9d40fffe;
    381: T0 = 32'h7fcf44b;
    382: T0 = 32'h2c8e57ff;
    383: T0 = 32'he076de54;
    384: T0 = 32'haa68343e;
    385: T0 = 32'h5a03ffe5;
    386: T0 = 32'h76e87b0f;
    387: T0 = 32'h46800fdf;
    388: T0 = 32'h7f7ff46;
    389: T0 = 32'h8d5cce0d;
    390: T0 = 32'hb07ba1aa;
    391: T0 = 32'h946bf37e;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T5 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T6 = reset ? 1'h0 : restartRegs_0;
  assign T7 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_11(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T5;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T6;
  reg  restartRegs_0;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (addr)
    0: T0 = 32'h9a277b02;
    1: T0 = 32'h487383e5;
    2: T0 = 32'hba85edc8;
    3: T0 = 32'h73c75718;
    4: T0 = 32'hb23ec5b3;
    5: T0 = 32'h3c05058c;
    6: T0 = 32'h3dc3f419;
    7: T0 = 32'h9940ff70;
    8: T0 = 32'h3fcd6627;
    9: T0 = 32'h71e205e1;
    10: T0 = 32'h53f83c20;
    11: T0 = 32'hf0fc01d0;
    12: T0 = 32'hf8ef80b1;
    13: T0 = 32'h8b5f001c;
    14: T0 = 32'he7ffc000;
    15: T0 = 32'hfe7da520;
    16: T0 = 32'h37e20080;
    17: T0 = 32'h61f4522;
    18: T0 = 32'h3b08000c;
    19: T0 = 32'h13dc;
    20: T0 = 32'h16420c0;
    21: T0 = 32'ha000013b;
    22: T0 = 32'h11b208;
    23: T0 = 32'hcf04401f;
    24: T0 = 32'h681fdb3;
    25: T0 = 32'h1d4077f3;
    26: T0 = 32'h1041ffa7;
    27: T0 = 32'h78a3f6ff;
    28: T0 = 32'hd201ffe3;
    29: T0 = 32'h3003677f;
    30: T0 = 32'hebf0fffc;
    31: T0 = 32'h8000e0ff;
    32: T0 = 32'h2bcffff;
    33: T0 = 32'hac008f4f;
    34: T0 = 32'h549ffe;
    35: T0 = 32'haff0c1f5;
    36: T0 = 32'hc00062ff;
    37: T0 = 32'h43ff8017;
    38: T0 = 32'hff8c3f3f;
    39: T0 = 32'hff8fc008;
    40: T0 = 32'hffff03f0;
    41: T0 = 32'hff089800;
    42: T0 = 32'h2fef0b0b;
    43: T0 = 32'hfffcdfd0;
    44: T0 = 32'hd1d7fff6;
    45: T0 = 32'hf7fdbc67;
    46: T0 = 32'hfd273f7f;
    47: T0 = 32'h681be9fe;
    48: T0 = 32'h173c5327;
    49: T0 = 32'h8998c54b;
    50: T0 = 32'h6fcfd3b5;
    51: T0 = 32'h9829931c;
    52: T0 = 32'h799817c5;
    53: T0 = 32'h6f6a5e04;
    54: T0 = 32'h47930059;
    55: T0 = 32'h1f602298;
    56: T0 = 32'h407f9030;
    57: T0 = 32'hfd447a1b;
    58: T0 = 32'h8e0141e5;
    59: T0 = 32'h3f920abe;
    60: T0 = 32'hfcc0ffc5;
    61: T0 = 32'h81e3b849;
    62: T0 = 32'hbf8303fe;
    63: T0 = 32'h740fc74b;
    64: T0 = 32'hfcf0d00f;
    65: T0 = 32'h4f804070;
    66: T0 = 32'h7a1e700;
    67: T0 = 32'h237c0007;
    68: T0 = 32'ha03e7e41;
    69: T0 = 32'h836f1e00;
    70: T0 = 32'h600303c1;
    71: T0 = 32'h38027bf8;
    72: T0 = 32'hb600807e;
    73: T0 = 32'h7fc0f63f;
    74: T0 = 32'h6a0fc0f;
    75: T0 = 32'h1ffcfff5;
    76: T0 = 32'hc0db7265;
    77: T0 = 32'hb27f7fc0;
    78: T0 = 32'hfc1e8b98;
    79: T0 = 32'hc52743f8;
    80: T0 = 32'h3dc726b9;
    81: T0 = 32'hfe19e43f;
    82: T0 = 32'hd3c8e497;
    83: T0 = 32'h1fed1d03;
    84: T0 = 32'h9e3e3c9a;
    85: T0 = 32'hc3f871ee;
    86: T0 = 32'ha8dbc3ce;
    87: T0 = 32'h3e077ebf;
    88: T0 = 32'h1b4ff036;
    89: T0 = 32'hcbe1766a;
    90: T0 = 32'h107fef81;
    91: T0 = 32'hec7e01d4;
    92: T0 = 32'he00a6370;
    93: T0 = 32'h328f4200;
    94: T0 = 32'h3e00e1bc;
    95: T0 = 32'hc9c0ea1;
    96: T0 = 32'ha2c03729;
    97: T0 = 32'h106f4a85;
    98: T0 = 32'hbc56bb7a;
    99: T0 = 32'h263bdc61;
    100: T0 = 32'h37635e31;
    101: T0 = 32'h8faa1012;
    102: T0 = 32'h7dfc28c1;
    103: T0 = 32'h7f8673;
    104: T0 = 32'h373ff611;
    105: T0 = 32'h2ffd3cd0;
    106: T0 = 32'hdbec4b90;
    107: T0 = 32'h6e1023ff;
    108: T0 = 32'haa0bf330;
    109: T0 = 32'h12ff4fff;
    110: T0 = 32'hff7eff00;
    111: T0 = 32'hf0fd3fff;
    112: T0 = 32'h7df7fffd;
    113: T0 = 32'h1ffa05ff;
    114: T0 = 32'hcdfefa7f;
    115: T0 = 32'hfeb8f07f;
    116: T0 = 32'hb7bfff0b;
    117: T0 = 32'hfbfdfcd5;
    118: T0 = 32'hf9e71fe3;
    119: T0 = 32'hfe7f3ffc;
    120: T0 = 32'hfc8fc1fe;
    121: T0 = 32'h5387c3ff;
    122: T0 = 32'hdfe3eca5;
    123: T0 = 32'h23217fb8;
    124: T0 = 32'ha0f002e8;
    125: T0 = 32'h74d3f0;
    126: T0 = 32'hfc00000;
    127: T0 = 32'h2dc43e;
    128: T0 = 32'h98103001;
    129: T0 = 32'h80071290;
    130: T0 = 32'h21000600;
    131: T0 = 32'hc1e;
    132: T0 = 32'h343a8020;
    133: T0 = 32'h400060e9;
    134: T0 = 32'h6438040;
    135: T0 = 32'h260008bc;
    136: T0 = 32'h3e4c43c;
    137: T0 = 32'h4b81c0ff;
    138: T0 = 32'h7f2f885;
    139: T0 = 32'hf7dedebf;
    140: T0 = 32'hc07fff61;
    141: T0 = 32'hffb30edf;
    142: T0 = 32'h573fffd1;
    143: T0 = 32'h7e01f1a9;
    144: T0 = 32'h198ffc58;
    145: T0 = 32'ha800d021;
    146: T0 = 32'h263587b2;
    147: T0 = 32'h51d27b24;
    148: T0 = 32'hf896d60;
    149: T0 = 32'h66cb1111;
    150: T0 = 32'h47f7637;
    151: T0 = 32'h99de1fbc;
    152: T0 = 32'hf50ff7c9;
    153: T0 = 32'he5994000;
    154: T0 = 32'h39078879;
    155: T0 = 32'hef52b042;
    156: T0 = 32'h16200061;
    157: T0 = 32'hf43de380;
    158: T0 = 32'hce01010d;
    159: T0 = 32'h798b0774;
    160: T0 = 32'h76900077;
    161: T0 = 32'h58c9c79a;
    162: T0 = 32'hfdeedc00;
    163: T0 = 32'hc5ff7543;
    164: T0 = 32'hf7a62e81;
    165: T0 = 32'hbfbf3f1c;
    166: T0 = 32'hfe38eaf0;
    167: T0 = 32'h79303f0;
    168: T0 = 32'h7f818d90;
    169: T0 = 32'h709f7f;
    170: T0 = 32'hafe0f0c9;
    171: T0 = 32'h768c7;
    172: T0 = 32'hfbfaff8f;
    173: T0 = 32'h20007719;
    174: T0 = 32'h7fe4e7f8;
    175: T0 = 32'h20f887fc;
    176: T0 = 32'hfff8b23f;
    177: T0 = 32'h261ffc6f;
    178: T0 = 32'hfffef8e1;
    179: T0 = 32'hebe10fe1;
    180: T0 = 32'hefffdffb;
    181: T0 = 32'hf80af81f;
    182: T0 = 32'hf1b72c43;
    183: T0 = 32'h48100;
    184: T0 = 32'hea3f0033;
    185: T0 = 32'hf8002be0;
    186: T0 = 32'hde990000;
    187: T0 = 32'h5e300844;
    188: T0 = 32'he8347200;
    189: T0 = 32'h97ea008f;
    190: T0 = 32'h710aa260;
    191: T0 = 32'hb09e280e;
    192: T0 = 32'h4d1ae010;
    193: T0 = 32'h8affb957;
    194: T0 = 32'hb9dc3c6c;
    195: T0 = 32'h6076a26a;
    196: T0 = 32'h1ecda72d;
    197: T0 = 32'h29296d5e;
    198: T0 = 32'hbb3ce35f;
    199: T0 = 32'h56c177f1;
    200: T0 = 32'h9db9f736;
    201: T0 = 32'h57e7059b;
    202: T0 = 32'h8fdeae00;
    203: T0 = 32'h1e3f21bc;
    204: T0 = 32'hff1bafc0;
    205: T0 = 32'h8181010e;
    206: T0 = 32'h3f1ff7bc;
    207: T0 = 32'he100fc07;
    208: T0 = 32'hf317a7;
    209: T0 = 32'h1b54bfe0;
    210: T0 = 32'h680ff;
    211: T0 = 32'hf1fdf9ff;
    212: T0 = 32'ha7f0fe06;
    213: T0 = 32'hce0f0c9f;
    214: T0 = 32'hfa3ffbf0;
    215: T0 = 32'hfee0c0d1;
    216: T0 = 32'h7f671f;
    217: T0 = 32'hbf86fe04;
    218: T0 = 32'h700ef834;
    219: T0 = 32'h1fc06ff9;
    220: T0 = 32'h380ee62;
    221: T0 = 32'h1f82af3;
    222: T0 = 32'h84fc3f40;
    223: T0 = 32'he0634177;
    224: T0 = 32'h7c0fe3fc;
    225: T0 = 32'hf7d0e019;
    226: T0 = 32'h5ffe9e1f;
    227: T0 = 32'hbffff807;
    228: T0 = 32'hfd9f2dc1;
    229: T0 = 32'hffff0f98;
    230: T0 = 32'hffd20354;
    231: T0 = 32'hfff01f2;
    232: T0 = 32'hfffb8500;
    233: T0 = 32'hfa3fa80d;
    234: T0 = 32'hff7dd280;
    235: T0 = 32'h9dc0084b;
    236: T0 = 32'hcfe2bf50;
    237: T0 = 32'he5f07067;
    238: T0 = 32'h97f3fde;
    239: T0 = 32'he0186001;
    240: T0 = 32'hd07503fd;
    241: T0 = 32'ha000f068;
    242: T0 = 32'h105c403f;
    243: T0 = 32'h67b89d4e;
    244: T0 = 32'h43c4a8db;
    245: T0 = 32'h118a7bdb;
    246: T0 = 32'h27ebccd1;
    247: T0 = 32'h4ffc51b4;
    248: T0 = 32'h911df20;
    249: T0 = 32'h98b08102;
    250: T0 = 32'hfffd4785;
    251: T0 = 32'hf3ad2280;
    252: T0 = 32'h5fff0015;
    253: T0 = 32'h3d3870;
    254: T0 = 32'h807f0001;
    255: T0 = 32'hed00e544;
    256: T0 = 32'h3030001;
    257: T0 = 32'h7fcfcf4;
    258: T0 = 32'hf8000133;
    259: T0 = 32'h807f1b62;
    260: T0 = 32'hffe0f880;
    261: T0 = 32'h480307a3;
    262: T0 = 32'h1fff86c0;
    263: T0 = 32'hf60c0fbf;
    264: T0 = 32'hd8fffeb8;
    265: T0 = 32'hfff0a3f9;
    266: T0 = 32'h6f6f8ccc;
    267: T0 = 32'hfff0e41f;
    268: T0 = 32'h67fff859;
    269: T0 = 32'hfc0fee63;
    270: T0 = 32'h163f7f87;
    271: T0 = 32'hff8056cd;
    272: T0 = 32'hbbbf8;
    273: T0 = 32'ha7c085e7;
    274: T0 = 32'h8016e31f;
    275: T0 = 32'h71407fbc;
    276: T0 = 32'h401702;
    277: T0 = 32'h43e01fb;
    278: T0 = 32'h801b00ac;
    279: T0 = 32'he0104004;
    280: T0 = 32'h53c70004;
    281: T0 = 32'hfc119000;
    282: T0 = 32'h92f40000;
    283: T0 = 32'h6fee0180;
    284: T0 = 32'hf8dc0000;
    285: T0 = 32'h51ff3fe6;
    286: T0 = 32'hff6e2300;
    287: T0 = 32'hf3f70fff;
    288: T0 = 32'h8fd727f0;
    289: T0 = 32'hee82cdff;
    290: T0 = 32'hffec9667;
    291: T0 = 32'h126a842;
    292: T0 = 32'h3fffacb3;
    293: T0 = 32'h48b07302;
    294: T0 = 32'h9a8f77f7;
    295: T0 = 32'h556bc76d;
    296: T0 = 32'h62bd7499;
    297: T0 = 32'hf67260c3;
    298: T0 = 32'h5d447000;
    299: T0 = 32'h60258e13;
    300: T0 = 32'h65284e40;
    301: T0 = 32'ha9d00956;
    302: T0 = 32'h458e0f0;
    303: T0 = 32'h2b8531af;
    304: T0 = 32'h1b3ba;
    305: T0 = 32'h8440fe04;
    306: T0 = 32'h70d1f83;
    307: T0 = 32'hf8e8fff0;
    308: T0 = 32'ha37d82b3;
    309: T0 = 32'h8f5187ff;
    310: T0 = 32'he817fe07;
    311: T0 = 32'hb87d964f;
    312: T0 = 32'h19802df0;
    313: T0 = 32'h78000d4;
    314: T0 = 32'h3c2007;
    315: T0 = 32'hc1bc780f;
    316: T0 = 32'he0464200;
    317: T0 = 32'hbf5fff80;
    318: T0 = 32'hffdc0ec0;
    319: T0 = 32'h881112fc;
    320: T0 = 32'h7ffff0a0;
    321: T0 = 32'hf025b27f;
    322: T0 = 32'h40fff5d3;
    323: T0 = 32'hfc0d3297;
    324: T0 = 32'h38033f6d;
    325: T0 = 32'h5800b74c;
    326: T0 = 32'h16091f4;
    327: T0 = 32'h400170f;
    328: T0 = 32'hec2ecf;
    329: T0 = 32'h40087efe;
    330: T0 = 32'h3951a8;
    331: T0 = 32'h1a7dd;
    332: T0 = 32'h4047a6fa;
    333: T0 = 32'hfc701e3f;
    334: T0 = 32'h10bfa30;
    335: T0 = 32'hbf1cc1e1;
    336: T0 = 32'h70011fcd;
    337: T0 = 32'h6fc4581;
    338: T0 = 32'h694001ff;
    339: T0 = 32'he57ee8f8;
    340: T0 = 32'h2648803f;
    341: T0 = 32'h9fe15fb4;
    342: T0 = 32'h940c5e62;
    343: T0 = 32'he029c3c8;
    344: T0 = 32'h57ce14b2;
    345: T0 = 32'h53c4adf;
    346: T0 = 32'h471e9f4c;
    347: T0 = 32'he89281ce;
    348: T0 = 32'h71bafda4;
    349: T0 = 32'h801c810f;
    350: T0 = 32'h100ffda;
    351: T0 = 32'h12bcc07;
    352: T0 = 32'h6c601ff8;
    353: T0 = 32'h42ac00;
    354: T0 = 32'h7683007f;
    355: T0 = 32'h6009f9e2;
    356: T0 = 32'h6ea44e2b;
    357: T0 = 32'h78018fc4;
    358: T0 = 32'h29d57ff;
    359: T0 = 32'hc16cf87f;
    360: T0 = 32'he0a8ebff;
    361: T0 = 32'hd97fff83;
    362: T0 = 32'hf4003fdf;
    363: T0 = 32'h6977ff0;
    364: T0 = 32'hfe0003f3;
    365: T0 = 32'h7c4247fc;
    366: T0 = 32'hc00c01f;
    367: T0 = 32'hfffeefe;
    368: T0 = 32'hec00ff11;
    369: T0 = 32'h1ff3ff3;
    370: T0 = 32'hfe583ce1;
    371: T0 = 32'h805f17c9;
    372: T0 = 32'hfe0007f7;
    373: T0 = 32'h22007238;
    374: T0 = 32'h2e009bff;
    375: T0 = 32'h4a6f327;
    376: T0 = 32'h52003a81;
    377: T0 = 32'h2e1f7a;
    378: T0 = 32'h7d830cb;
    379: T0 = 32'h861ff;
    380: T0 = 32'hc8ed918f;
    381: T0 = 32'h4881f1b7;
    382: T0 = 32'hf98d7dbe;
    383: T0 = 32'h4f3f3ba8;
    384: T0 = 32'h7fcb6d9a;
    385: T0 = 32'h77cddfbb;
    386: T0 = 32'h5ff39bdd;
    387: T0 = 32'hbbd6fb7e;
    388: T0 = 32'h4cf2ec23;
    389: T0 = 32'he66b99bc;
    390: T0 = 32'ha10523c;
    391: T0 = 32'hf19822bb;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T5 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T6 = reset ? 1'h0 : restartRegs_0;
  assign T7 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_12(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T5;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T6;
  reg  restartRegs_0;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (addr)
    0: T0 = 32'hef8f5d53;
    1: T0 = 32'hc7f0d52f;
    2: T0 = 32'hd7b0e727;
    3: T0 = 32'h9c1c529a;
    4: T0 = 32'h1ca88ccb;
    5: T0 = 32'hc202001b;
    6: T0 = 32'h12a3f5fc;
    7: T0 = 32'heb00c07d;
    8: T0 = 32'h1047cd3f;
    9: T0 = 32'h43f9ca02;
    10: T0 = 32'hff430167;
    11: T0 = 32'hd2f7c12;
    12: T0 = 32'hff847c22;
    13: T0 = 32'h8d6fc1;
    14: T0 = 32'h7ff01fc7;
    15: T0 = 32'h3084727c;
    16: T0 = 32'h85e6e1fa;
    17: T0 = 32'h1c0fb8f;
    18: T0 = 32'h81c0ff01;
    19: T0 = 32'h1f06d0;
    20: T0 = 32'hfc3057f0;
    21: T0 = 32'h3c01e;
    22: T0 = 32'hffe3afff;
    23: T0 = 32'h180cdf00;
    24: T0 = 32'hffbe1adf;
    25: T0 = 32'hc5f17ff8;
    26: T0 = 32'hff9c13e;
    27: T0 = 32'hf817c01f;
    28: T0 = 32'ha03ffe0f;
    29: T0 = 32'hff8ac400;
    30: T0 = 32'hc2830ff1;
    31: T0 = 32'hff91fc0;
    32: T0 = 32'h84b8003e;
    33: T0 = 32'h807fff24;
    34: T0 = 32'hf23dd030;
    35: T0 = 32'h1d008ffd;
    36: T0 = 32'h80f0dbcc;
    37: T0 = 32'ha5fc82ff;
    38: T0 = 32'hf000e4df;
    39: T0 = 32'h3afd871;
    40: T0 = 32'hff589dc8;
    41: T0 = 32'h80afe81f;
    42: T0 = 32'hfc8f877;
    43: T0 = 32'h1007e7cf;
    44: T0 = 32'he7fd7803;
    45: T0 = 32'hc20084f0;
    46: T0 = 32'h6dad3a46;
    47: T0 = 32'h280221f9;
    48: T0 = 32'h833ff5a9;
    49: T0 = 32'hf110c07c;
    50: T0 = 32'h125e4c4c;
    51: T0 = 32'ha61b3dbf;
    52: T0 = 32'hd3ec4524;
    53: T0 = 32'hf5fe3a0a;
    54: T0 = 32'haf347cf9;
    55: T0 = 32'hfe8daff0;
    56: T0 = 32'h43705de;
    57: T0 = 32'h1ec2307c;
    58: T0 = 32'h9403c060;
    59: T0 = 32'hfff68d3f;
    60: T0 = 32'he6cafe1c;
    61: T0 = 32'hc0ffb02d;
    62: T0 = 32'hfa416de1;
    63: T0 = 32'h80031d80;
    64: T0 = 32'hfff8a7e;
    65: T0 = 32'hda00f0fd;
    66: T0 = 32'h7ffe67;
    67: T0 = 32'hfe803f87;
    68: T0 = 32'h170798;
    69: T0 = 32'hffec63f8;
    70: T0 = 32'hc401c03e;
    71: T0 = 32'h1eff9e7f;
    72: T0 = 32'he5f9fc03;
    73: T0 = 32'hf1ffe287;
    74: T0 = 32'hf83f7fe3;
    75: T0 = 32'hff9ecc6c;
    76: T0 = 32'he07b43ee;
    77: T0 = 32'h9ff9c01c;
    78: T0 = 32'hdfe7603e;
    79: T0 = 32'hc1fbc801;
    80: T0 = 32'h8bf31de0;
    81: T0 = 32'h85df0200;
    82: T0 = 32'hf83f0390;
    83: T0 = 32'hfe74e028;
    84: T0 = 32'h5fc1c02a;
    85: T0 = 32'h79739800;
    86: T0 = 32'h3d7c00cb;
    87: T0 = 32'he23b3ea1;
    88: T0 = 32'hb8b3200b;
    89: T0 = 32'hff330108;
    90: T0 = 32'hd7b73008;
    91: T0 = 32'h8ffc04ef;
    92: T0 = 32'ha8172020;
    93: T0 = 32'hb47f03ff;
    94: T0 = 32'he000fc83;
    95: T0 = 32'h63ef63bf;
    96: T0 = 32'h7e00a70f;
    97: T0 = 32'h8c22feb5;
    98: T0 = 32'ha6bda3e7;
    99: T0 = 32'h7f49b8b2;
    100: T0 = 32'hf472b1ec;
    101: T0 = 32'hf7405e46;
    102: T0 = 32'h650b6883;
    103: T0 = 32'hb7e94363;
    104: T0 = 32'hc2a5e05f;
    105: T0 = 32'h1effff9c;
    106: T0 = 32'hff1603d8;
    107: T0 = 32'hebdff887;
    108: T0 = 32'hffff6541;
    109: T0 = 32'he9a90000;
    110: T0 = 32'h7fff03c7;
    111: T0 = 32'hffba7400;
    112: T0 = 32'h71ff007f;
    113: T0 = 32'hfffb7f10;
    114: T0 = 32'h52190001;
    115: T0 = 32'h7d4fc5;
    116: T0 = 32'hcb461602;
    117: T0 = 32'h74011202;
    118: T0 = 32'hf504010;
    119: T0 = 32'h67801e82;
    120: T0 = 32'h307a0001;
    121: T0 = 32'hb8f811fe;
    122: T0 = 32'h8387e698;
    123: T0 = 32'h7edfef3f;
    124: T0 = 32'hf8b8fe09;
    125: T0 = 32'hc720b2f3;
    126: T0 = 32'h83c6dfbc;
    127: T0 = 32'h7ef8a3ff;
    128: T0 = 32'hcf3cfcaf;
    129: T0 = 32'he1fef97d;
    130: T0 = 32'hfe0fffdf;
    131: T0 = 32'h7f8fffaf;
    132: T0 = 32'hff53ffff;
    133: T0 = 32'h53f1fffc;
    134: T0 = 32'hfffeb3ff;
    135: T0 = 32'h833f97ef;
    136: T0 = 32'hffff75de;
    137: T0 = 32'hec138000;
    138: T0 = 32'hf1fd01eb;
    139: T0 = 32'h80b07000;
    140: T0 = 32'he71f0030;
    141: T0 = 32'hfe549950;
    142: T0 = 32'h6d03000e;
    143: T0 = 32'hffe63d65;
    144: T0 = 32'h4e3a013;
    145: T0 = 32'h247d46a6;
    146: T0 = 32'h7b115379;
    147: T0 = 32'haaff845f;
    148: T0 = 32'h780660fb;
    149: T0 = 32'he81760d;
    150: T0 = 32'hf49fa5c7;
    151: T0 = 32'hb0924ffe;
    152: T0 = 32'h97fdf816;
    153: T0 = 32'he5e21fff;
    154: T0 = 32'ha37ffff7;
    155: T0 = 32'hefef1dff;
    156: T0 = 32'h2136fffc;
    157: T0 = 32'h60f1f9af;
    158: T0 = 32'h1b801fff;
    159: T0 = 32'h1dff879;
    160: T0 = 32'hc548201f;
    161: T0 = 32'hbf1cb0;
    162: T0 = 32'hcd0d9c00;
    163: T0 = 32'hc;
    164: T0 = 32'h1f06940;
    165: T0 = 32'he0001001;
    166: T0 = 32'h30320;
    167: T0 = 32'h1330e586;
    168: T0 = 32'hb3fce00a;
    169: T0 = 32'hfc12b7b7;
    170: T0 = 32'h331f7e08;
    171: T0 = 32'hffc1689c;
    172: T0 = 32'hdbee0e0;
    173: T0 = 32'hf7fe349c;
    174: T0 = 32'h1c75f0f;
    175: T0 = 32'hf7bf7427;
    176: T0 = 32'h80119008;
    177: T0 = 32'h87ff03d3;
    178: T0 = 32'hf0079e9b;
    179: T0 = 32'hf87bff1e;
    180: T0 = 32'hff00f8a7;
    181: T0 = 32'h1fa55cff;
    182: T0 = 32'h6de0ff8f;
    183: T0 = 32'hf7e7eff;
    184: T0 = 32'he3e8ffff;
    185: T0 = 32'h16ef00d;
    186: T0 = 32'hc45dbfff;
    187: T0 = 32'hf0147f00;
    188: T0 = 32'h57ff26bf;
    189: T0 = 32'h9600f3ff;
    190: T0 = 32'h1f9de10f;
    191: T0 = 32'h4f0f0fd;
    192: T0 = 32'ha7f9c719;
    193: T0 = 32'ha3eec401;
    194: T0 = 32'h71ef17d8;
    195: T0 = 32'he495459;
    196: T0 = 32'h12a4b2a2;
    197: T0 = 32'ha498eb4b;
    198: T0 = 32'h2b0d0a1f;
    199: T0 = 32'h6a9cf3b8;
    200: T0 = 32'h8aba2a5;
    201: T0 = 32'h15100667;
    202: T0 = 32'hd45f3133;
    203: T0 = 32'h2021e4fb;
    204: T0 = 32'h502a2923;
    205: T0 = 32'h7d01199b;
    206: T0 = 32'h1f8dc678;
    207: T0 = 32'hd69f1cd;
    208: T0 = 32'h9b881ecf;
    209: T0 = 32'h263790c;
    210: T0 = 32'h389cf5ff;
    211: T0 = 32'h28035f80;
    212: T0 = 32'h4fe9079a;
    213: T0 = 32'h838013fe;
    214: T0 = 32'ha3d01ff;
    215: T0 = 32'hf81be3ef;
    216: T0 = 32'hf067e17f;
    217: T0 = 32'hff87fe1d;
    218: T0 = 32'hff05bc07;
    219: T0 = 32'hdbe37fc1;
    220: T0 = 32'h1ff015c0;
    221: T0 = 32'h69c03f8;
    222: T0 = 32'h83ff81ec;
    223: T0 = 32'he0538219;
    224: T0 = 32'ha83f801f;
    225: T0 = 32'hf800e081;
    226: T0 = 32'h2f830c07;
    227: T0 = 32'h7780fe12;
    228: T0 = 32'ha020e0;
    229: T0 = 32'h7c00789;
    230: T0 = 32'hf47c14f;
    231: T0 = 32'ha07cf0f8;
    232: T0 = 32'hc1ffe000;
    233: T0 = 32'hd7077f03;
    234: T0 = 32'h322ecfc4;
    235: T0 = 32'h91385ff0;
    236: T0 = 32'h3fd9134;
    237: T0 = 32'h91a0ceff;
    238: T0 = 32'h303ff0ca;
    239: T0 = 32'hbea8538f;
    240: T0 = 32'hbe07ff49;
    241: T0 = 32'he0611848;
    242: T0 = 32'h36306ebe;
    243: T0 = 32'h4e087425;
    244: T0 = 32'h5f2fcf47;
    245: T0 = 32'h57cbffc5;
    246: T0 = 32'hef776ace;
    247: T0 = 32'hc3ee3df3;
    248: T0 = 32'h82b0b3c3;
    249: T0 = 32'hed9c483e;
    250: T0 = 32'hc172f6cf;
    251: T0 = 32'he033100b;
    252: T0 = 32'hd3ff02bd;
    253: T0 = 32'h77ef1780;
    254: T0 = 32'h4bb90001;
    255: T0 = 32'hfc6936be;
    256: T0 = 32'hf167fc00;
    257: T0 = 32'h45c10337;
    258: T0 = 32'h90589ffe;
    259: T0 = 32'hc01f837;
    260: T0 = 32'h1defb7ff;
    261: T0 = 32'h7580cfc1;
    262: T0 = 32'hf02008ff;
    263: T0 = 32'hfff887e;
    264: T0 = 32'hfff2f07f;
    265: T0 = 32'hf8e3600f;
    266: T0 = 32'h3fffef03;
    267: T0 = 32'h9e03da00;
    268: T0 = 32'h33ff1e78;
    269: T0 = 32'ha0018360;
    270: T0 = 32'h1fdf01e3;
    271: T0 = 32'hfa0000f3;
    272: T0 = 32'h7ff700e;
    273: T0 = 32'h37f86007;
    274: T0 = 32'h83fb6400;
    275: T0 = 32'hdc007c0;
    276: T0 = 32'h27ff8ad0;
    277: T0 = 32'hff3c0264;
    278: T0 = 32'hc87f681f;
    279: T0 = 32'hffa58006;
    280: T0 = 32'h3a172f03;
    281: T0 = 32'hffe66207;
    282: T0 = 32'h35804040;
    283: T0 = 32'h30f49300;
    284: T0 = 32'h67e1612;
    285: T0 = 32'h40f0ce5a;
    286: T0 = 32'h746097;
    287: T0 = 32'h64e08029;
    288: T0 = 32'h90196906;
    289: T0 = 32'h7445f85c;
    290: T0 = 32'h27508;
    291: T0 = 32'h399003f8;
    292: T0 = 32'h194a1;
    293: T0 = 32'h1db3648d;
    294: T0 = 32'h4191c67a;
    295: T0 = 32'hebd4a05;
    296: T0 = 32'h89277725;
    297: T0 = 32'heb20a91f;
    298: T0 = 32'h84b81889;
    299: T0 = 32'h7b11884;
    300: T0 = 32'h395d0000;
    301: T0 = 32'h7ffe2031;
    302: T0 = 32'h6fac6600;
    303: T0 = 32'hf3757ea2;
    304: T0 = 32'h5010301;
    305: T0 = 32'h10045200;
    306: T0 = 32'h47e00038;
    307: T0 = 32'hf80e00;
    308: T0 = 32'hc0180004;
    309: T0 = 32'ha2dfc;
    310: T0 = 32'hc000fb81;
    311: T0 = 32'h95bf;
    312: T0 = 32'h9e7cffff;
    313: T0 = 32'hfc02ff58;
    314: T0 = 32'hff6703df;
    315: T0 = 32'h3fffffff;
    316: T0 = 32'hfff9901e;
    317: T0 = 32'heeff7ebf;
    318: T0 = 32'h9fffe520;
    319: T0 = 32'hfb6f07e1;
    320: T0 = 32'h4bff1386;
    321: T0 = 32'hffacd03f;
    322: T0 = 32'hc07ff73c;
    323: T0 = 32'hff745281;
    324: T0 = 32'h30ff5;
    325: T0 = 32'h1ff86a48;
    326: T0 = 32'hebc0807f;
    327: T0 = 32'hff2c6a;
    328: T0 = 32'hfd98e800;
    329: T0 = 32'h93b10006;
    330: T0 = 32'h1e3ff0;
    331: T0 = 32'haedce000;
    332: T0 = 32'h9800069f;
    333: T0 = 32'h1313ff60;
    334: T0 = 32'h3860cbb2;
    335: T0 = 32'hb0270fff;
    336: T0 = 32'h67c00002;
    337: T0 = 32'hac0aefbe;
    338: T0 = 32'h96fb0204;
    339: T0 = 32'hb8403ada;
    340: T0 = 32'h69dec77e;
    341: T0 = 32'ha62a46ae;
    342: T0 = 32'hac25235f;
    343: T0 = 32'he5088258;
    344: T0 = 32'h5beb6c53;
    345: T0 = 32'hbb808d1d;
    346: T0 = 32'hd4c51115;
    347: T0 = 32'he52c7f80;
    348: T0 = 32'hec100d43;
    349: T0 = 32'he8481df8;
    350: T0 = 32'h7fc9801d;
    351: T0 = 32'hbcd1eb6b;
    352: T0 = 32'hc27efc09;
    353: T0 = 32'hf9f836be;
    354: T0 = 32'ha681c7c0;
    355: T0 = 32'hf144661;
    356: T0 = 32'hf86a3f39;
    357: T0 = 32'he039c0e4;
    358: T0 = 32'hf843fd3;
    359: T0 = 32'h86001f0d;
    360: T0 = 32'hfc1938;
    361: T0 = 32'hf6c080ff;
    362: T0 = 32'hfd4ab;
    363: T0 = 32'hffd5f007;
    364: T0 = 32'h37783ffa;
    365: T0 = 32'hfe89600;
    366: T0 = 32'h5aff01fe;
    367: T0 = 32'hf07fec00;
    368: T0 = 32'hf38f4007;
    369: T0 = 32'hff072fdf;
    370: T0 = 32'h7bc80c40;
    371: T0 = 32'h26600087;
    372: T0 = 32'h7a44de4;
    373: T0 = 32'h51734008;
    374: T0 = 32'hf87df28f;
    375: T0 = 32'h1c017f00;
    376: T0 = 32'h3b871c6c;
    377: T0 = 32'h30de47e8;
    378: T0 = 32'hb0987fce;
    379: T0 = 32'hc011aef7;
    380: T0 = 32'h930dcfe2;
    381: T0 = 32'h9c03015b;
    382: T0 = 32'h3ab37ff8;
    383: T0 = 32'h73e0e000;
    384: T0 = 32'h180079a;
    385: T0 = 32'h2a3ef73c;
    386: T0 = 32'hc038a6c5;
    387: T0 = 32'h9d3ffffb;
    388: T0 = 32'hfd04ac17;
    389: T0 = 32'he3357f7e;
    390: T0 = 32'h1fbebd0b;
    391: T0 = 32'haeb9cc5e;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T5 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T6 = reset ? 1'h0 : restartRegs_0;
  assign T7 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_13(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T5;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T6;
  reg  restartRegs_0;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (addr)
    0: T0 = 32'he5fbce98;
    1: T0 = 32'hc5cd10d2;
    2: T0 = 32'hedd2d6e1;
    3: T0 = 32'h1c0097d9;
    4: T0 = 32'he99dc2a;
    5: T0 = 32'hc004fbc3;
    6: T0 = 32'h9950bc0;
    7: T0 = 32'h20005f8c;
    8: T0 = 32'h1589e;
    9: T0 = 32'h1d00f170;
    10: T0 = 32'h38da0;
    11: T0 = 32'h70a80f09;
    12: T0 = 32'hc0007c43;
    13: T0 = 32'h25d723e0;
    14: T0 = 32'h7c0007ad;
    15: T0 = 32'h31f588ff;
    16: T0 = 32'h8ffdf828;
    17: T0 = 32'hfff3ac97;
    18: T0 = 32'ha53eff82;
    19: T0 = 32'hffff0369;
    20: T0 = 32'hff0f7ffc;
    21: T0 = 32'h60fbf01a;
    22: T0 = 32'h9ffffb71;
    23: T0 = 32'hc0f0f80;
    24: T0 = 32'h71ff0071;
    25: T0 = 32'hd06032fe;
    26: T0 = 32'h471fa0b7;
    27: T0 = 32'h6ce2d05f;
    28: T0 = 32'hc270fc00;
    29: T0 = 32'h93e1a789;
    30: T0 = 32'hf6071fdf;
    31: T0 = 32'h3dbc57d0;
    32: T0 = 32'hdd09c078;
    33: T0 = 32'h80c1f16b;
    34: T0 = 32'h10d0b43;
    35: T0 = 32'hc0003ef3;
    36: T0 = 32'h6beb4;
    37: T0 = 32'h582001e7;
    38: T0 = 32'heb3c;
    39: T0 = 32'h6f6a41f;
    40: T0 = 32'hd000ff7a;
    41: T0 = 32'h40674200;
    42: T0 = 32'hbf0183f8;
    43: T0 = 32'ha1d7001;
    44: T0 = 32'h7170007e;
    45: T0 = 32'he70144c0;
    46: T0 = 32'hc1fc820a;
    47: T0 = 32'heaee2cef;
    48: T0 = 32'hec8e6a96;
    49: T0 = 32'h180108c2;
    50: T0 = 32'h751a7d91;
    51: T0 = 32'hc598a04;
    52: T0 = 32'ha0bb022a;
    53: T0 = 32'hb7867ee4;
    54: T0 = 32'h5e01bd7a;
    55: T0 = 32'h58a5c17f;
    56: T0 = 32'h3900fc9e;
    57: T0 = 32'he1bac12;
    58: T0 = 32'hb60027e2;
    59: T0 = 32'he7888543;
    60: T0 = 32'he8f1fff;
    61: T0 = 32'hfcfcf047;
    62: T0 = 32'ha08fa54f;
    63: T0 = 32'h5f9f3c07;
    64: T0 = 32'hf807c580;
    65: T0 = 32'h23fc03c1;
    66: T0 = 32'hc7c0014c;
    67: T0 = 32'hfdff001c;
    68: T0 = 32'hfc7dc23c;
    69: T0 = 32'hffdf0081;
    70: T0 = 32'h3fc70c01;
    71: T0 = 32'h7ff009df;
    72: T0 = 32'h6a3cfbc0;
    73: T0 = 32'hc77f01f9;
    74: T0 = 32'hf1610ffc;
    75: T0 = 32'h663e1be;
    76: T0 = 32'h3b445ff;
    77: T0 = 32'h8052fe03;
    78: T0 = 32'h1e1cdf;
    79: T0 = 32'hbc01fbf0;
    80: T0 = 32'h380307f3;
    81: T0 = 32'h7a686f8f;
    82: T0 = 32'h8665ed;
    83: T0 = 32'h6f979afc;
    84: T0 = 32'haff0c0fe;
    85: T0 = 32'h5f8d77f;
    86: T0 = 32'hf97dfeab;
    87: T0 = 32'he00f1e49;
    88: T0 = 32'hfe1f1f9c;
    89: T0 = 32'hff3e011a;
    90: T0 = 32'he7ea03f2;
    91: T0 = 32'h9dff3700;
    92: T0 = 32'h4267e6bc;
    93: T0 = 32'hda7e414a;
    94: T0 = 32'hef726f4b;
    95: T0 = 32'hd56f1040;
    96: T0 = 32'h6e094058;
    97: T0 = 32'h1bc4e2d1;
    98: T0 = 32'h518ec1c4;
    99: T0 = 32'h95142e55;
    100: T0 = 32'h2c234063;
    101: T0 = 32'h1e18cb6a;
    102: T0 = 32'h9e03e26;
    103: T0 = 32'h9175190e;
    104: T0 = 32'hfd73efe0;
    105: T0 = 32'h8017006d;
    106: T0 = 32'hfeeba7fb;
    107: T0 = 32'he6092007;
    108: T0 = 32'hdbf5feff;
    109: T0 = 32'h9241e001;
    110: T0 = 32'h53f9f81;
    111: T0 = 32'hf884fc00;
    112: T0 = 32'h84041f79;
    113: T0 = 32'h87c78f00;
    114: T0 = 32'h7e5001f2;
    115: T0 = 32'hfc3e81a0;
    116: T0 = 32'hf16f003f;
    117: T0 = 32'h7fc3f9e6;
    118: T0 = 32'h1fdbc037;
    119: T0 = 32'hdbf83fcc;
    120: T0 = 32'hc1f44c07;
    121: T0 = 32'h9781e9fc;
    122: T0 = 32'h440f8247;
    123: T0 = 32'hf8fc7e1f;
    124: T0 = 32'hcc40f0c6;
    125: T0 = 32'hfb30ff9;
    126: T0 = 32'h7ce6df01;
    127: T0 = 32'h62f66cfe;
    128: T0 = 32'h77cfe3c0;
    129: T0 = 32'h6617010b;
    130: T0 = 32'hb9bf2f3c;
    131: T0 = 32'hfc7383e0;
    132: T0 = 32'hcb30031;
    133: T0 = 32'hffc6103a;
    134: T0 = 32'he2be76fb;
    135: T0 = 32'hd3fd58c2;
    136: T0 = 32'hec1f2945;
    137: T0 = 32'h7d4743f4;
    138: T0 = 32'hff030346;
    139: T0 = 32'hefb0a5fe;
    140: T0 = 32'h8ffcf024;
    141: T0 = 32'hf6e99f;
    142: T0 = 32'hf2fefc06;
    143: T0 = 32'hc1530539;
    144: T0 = 32'h15af4fe3;
    145: T0 = 32'h7e018a00;
    146: T0 = 32'h1e98707c;
    147: T0 = 32'h3f3832bb;
    148: T0 = 32'ha7721769;
    149: T0 = 32'hb21dd957;
    150: T0 = 32'h50768761;
    151: T0 = 32'h5dd07fe;
    152: T0 = 32'h61822fa5;
    153: T0 = 32'h528df0fd;
    154: T0 = 32'h89c0844a;
    155: T0 = 32'h2f5603;
    156: T0 = 32'h2d66081b;
    157: T0 = 32'ha0083690;
    158: T0 = 32'h13de01e0;
    159: T0 = 32'hf000c330;
    160: T0 = 32'hffad001f;
    161: T0 = 32'h3e03f33d;
    162: T0 = 32'h3fffe800;
    163: T0 = 32'hbdc0070e;
    164: T0 = 32'h7ffd787;
    165: T0 = 32'hfe3c387b;
    166: T0 = 32'h807fff6c;
    167: T0 = 32'hff4777c7;
    168: T0 = 32'hd80fc7f1;
    169: T0 = 32'hf96915ff;
    170: T0 = 32'h6381fc7f;
    171: T0 = 32'h7fa5ea3f;
    172: T0 = 32'h1918ffc3;
    173: T0 = 32'hc1fa7f63;
    174: T0 = 32'he403e774;
    175: T0 = 32'hff4fc09c;
    176: T0 = 32'hfacb0a01;
    177: T0 = 32'h97f00e00;
    178: T0 = 32'h7f803a4;
    179: T0 = 32'hcebf4de0;
    180: T0 = 32'hfabf000c;
    181: T0 = 32'h87f01ef;
    182: T0 = 32'hbfd8f002;
    183: T0 = 32'h3a60f;
    184: T0 = 32'h78765e00;
    185: T0 = 32'h4cce08d0;
    186: T0 = 32'h46a8000;
    187: T0 = 32'h300562;
    188: T0 = 32'h6400c780;
    189: T0 = 32'h233501fe;
    190: T0 = 32'h411141ff;
    191: T0 = 32'hdaaff7f;
    192: T0 = 32'hf000e657;
    193: T0 = 32'h7b8226c1;
    194: T0 = 32'hbd44be81;
    195: T0 = 32'h2e14d48c;
    196: T0 = 32'h6af08505;
    197: T0 = 32'h9af491bd;
    198: T0 = 32'h11f9dce0;
    199: T0 = 32'h7b25e560;
    200: T0 = 32'he1a10100;
    201: T0 = 32'hc1fb36e3;
    202: T0 = 32'hee748000;
    203: T0 = 32'hc07f0133;
    204: T0 = 32'hff419c80;
    205: T0 = 32'h3c070003;
    206: T0 = 32'hde700725;
    207: T0 = 32'h9587e8f0;
    208: T0 = 32'hfcc1df;
    209: T0 = 32'he079ff7f;
    210: T0 = 32'h400ffc06;
    211: T0 = 32'h3c4a0fff;
    212: T0 = 32'h2200ffc0;
    213: T0 = 32'h1f0e33f;
    214: T0 = 32'hbe50fc3d;
    215: T0 = 32'hf00ffeab;
    216: T0 = 32'h7eed7fe3;
    217: T0 = 32'h1ff83ff2;
    218: T0 = 32'h87ffc6fe;
    219: T0 = 32'he9ffa1ff;
    220: T0 = 32'h807feb27;
    221: T0 = 32'hfe3e020f;
    222: T0 = 32'hf2075966;
    223: T0 = 32'h7f911000;
    224: T0 = 32'hf000019;
    225: T0 = 32'h2aaba00;
    226: T0 = 32'hee9800c2;
    227: T0 = 32'hc083c780;
    228: T0 = 32'hca0b004c;
    229: T0 = 32'h3c0d5c0c;
    230: T0 = 32'hd09bc056;
    231: T0 = 32'hae02143;
    232: T0 = 32'h814f3b84;
    233: T0 = 32'hdb2b0024;
    234: T0 = 32'h58164130;
    235: T0 = 32'hb87801f;
    236: T0 = 32'h6580e06b;
    237: T0 = 32'h7a83901;
    238: T0 = 32'h86bcf802;
    239: T0 = 32'hc16d34bf;
    240: T0 = 32'h7efffe00;
    241: T0 = 32'hfc075b5f;
    242: T0 = 32'h70c7bc62;
    243: T0 = 32'hdfc187fb;
    244: T0 = 32'h3ff26f58;
    245: T0 = 32'haea8278d;
    246: T0 = 32'h41dcae65;
    247: T0 = 32'ha27c57c1;
    248: T0 = 32'hdabf08b1;
    249: T0 = 32'hea1a84b9;
    250: T0 = 32'h814f9510;
    251: T0 = 32'hf333650c;
    252: T0 = 32'h501b3e19;
    253: T0 = 32'hbfc39f00;
    254: T0 = 32'hae0b01c8;
    255: T0 = 32'h39ff813e;
    256: T0 = 32'he7c1e80f;
    257: T0 = 32'h78ff81b;
    258: T0 = 32'h7facfe00;
    259: T0 = 32'h43fc0f83;
    260: T0 = 32'hc3e497fa;
    261: T0 = 32'hd80ff0f0;
    262: T0 = 32'hf83faa3f;
    263: T0 = 32'hf385ff0f;
    264: T0 = 32'h3783f807;
    265: T0 = 32'h3fa0fe31;
    266: T0 = 32'h87f81f6e;
    267: T0 = 32'h83f78690;
    268: T0 = 32'h77fb41ff;
    269: T0 = 32'h303fe01c;
    270: T0 = 32'hf4fef68f;
    271: T0 = 32'hc7a3742f;
    272: T0 = 32'h9fcb8804;
    273: T0 = 32'h7e5a4370;
    274: T0 = 32'ha4ee20a0;
    275: T0 = 32'h5bef061e;
    276: T0 = 32'hcc17e99f;
    277: T0 = 32'h2dff1873;
    278: T0 = 32'hf8c1843b;
    279: T0 = 32'hcab05c7;
    280: T0 = 32'h7f2c7802;
    281: T0 = 32'ha078f074;
    282: T0 = 32'hbf723c2;
    283: T0 = 32'hd077a945;
    284: T0 = 32'hf61f2be0;
    285: T0 = 32'hfe0000c2;
    286: T0 = 32'h2d20913f;
    287: T0 = 32'h8fe0f01a;
    288: T0 = 32'h1bbbc87;
    289: T0 = 32'hb4ff1c03;
    290: T0 = 32'h3ffda5b8;
    291: T0 = 32'hd1a43060;
    292: T0 = 32'h87f02aa;
    293: T0 = 32'h3631a018;
    294: T0 = 32'hd98b8f4a;
    295: T0 = 32'h4e5d4f9;
    296: T0 = 32'h639a6c78;
    297: T0 = 32'h9ddcab2a;
    298: T0 = 32'hacbd3790;
    299: T0 = 32'h9dfff7bd;
    300: T0 = 32'hb98a1dfd;
    301: T0 = 32'h90c102f0;
    302: T0 = 32'h2369f51e;
    303: T0 = 32'hf09e1f7;
    304: T0 = 32'hf12ee5f;
    305: T0 = 32'hc5c5f80f;
    306: T0 = 32'h66ffce;
    307: T0 = 32'h59a23f01;
    308: T0 = 32'hc00202f9;
    309: T0 = 32'h961e3ff4;
    310: T0 = 32'h77ef0003;
    311: T0 = 32'hff4700fe;
    312: T0 = 32'h677fe130;
    313: T0 = 32'hff1d80f7;
    314: T0 = 32'h3aa7fc17;
    315: T0 = 32'hbfc03f0c;
    316: T0 = 32'hdab3c0;
    317: T0 = 32'h97e001fd;
    318: T0 = 32'h7ef53c;
    319: T0 = 32'hec5ef10f;
    320: T0 = 32'hc80f3fd1;
    321: T0 = 32'hfec09f98;
    322: T0 = 32'he00380f2;
    323: T0 = 32'hffedfdfe;
    324: T0 = 32'h1a20fc0f;
    325: T0 = 32'h1ffaffc7;
    326: T0 = 32'h80703fc0;
    327: T0 = 32'h41ff0f5c;
    328: T0 = 32'he016f19e;
    329: T0 = 32'ha3fc17a;
    330: T0 = 32'h90162043;
    331: T0 = 32'h7a877c9f;
    332: T0 = 32'h7b442218;
    333: T0 = 32'he6e83fbb;
    334: T0 = 32'h86bf0052;
    335: T0 = 32'hb455c5a2;
    336: T0 = 32'ha06cad55;
    337: T0 = 32'hd017af59;
    338: T0 = 32'h8a0c1ba1;
    339: T0 = 32'he018b570;
    340: T0 = 32'h3aac0228;
    341: T0 = 32'h6f019d16;
    342: T0 = 32'h1ab4ef67;
    343: T0 = 32'h248ef95;
    344: T0 = 32'h44387ad;
    345: T0 = 32'hf5e52f3b;
    346: T0 = 32'hec3558ce;
    347: T0 = 32'hfc105eff;
    348: T0 = 32'he2aa71b7;
    349: T0 = 32'hf9889edf;
    350: T0 = 32'hd80fc2a9;
    351: T0 = 32'hb7c9ecdd;
    352: T0 = 32'he042807c;
    353: T0 = 32'hffffd567;
    354: T0 = 32'h7d40519f;
    355: T0 = 32'h9cf7ffc7;
    356: T0 = 32'hc20fb0ff;
    357: T0 = 32'hfa017ffe;
    358: T0 = 32'h3a45cdf8;
    359: T0 = 32'h63f80041;
    360: T0 = 32'ha3c40504;
    361: T0 = 32'hfd1f0000;
    362: T0 = 32'hfc3f0076;
    363: T0 = 32'hfe471418;
    364: T0 = 32'hffc3e004;
    365: T0 = 32'h7fb9f81;
    366: T0 = 32'he5e8bf80;
    367: T0 = 32'h1ffa55;
    368: T0 = 32'hf83e1fff;
    369: T0 = 32'he040ffe4;
    370: T0 = 32'hf6fa4ff;
    371: T0 = 32'h3f06ffea;
    372: T0 = 32'h61ff4603;
    373: T0 = 32'hf7f00ffe;
    374: T0 = 32'h85ff811c;
    375: T0 = 32'hf6bf707f;
    376: T0 = 32'hfc7f0252;
    377: T0 = 32'hff7b4bf0;
    378: T0 = 32'hffcf8008;
    379: T0 = 32'h9fc74cff;
    380: T0 = 32'h71ffc000;
    381: T0 = 32'hfc7808df;
    382: T0 = 32'h3115000;
    383: T0 = 32'hde785094;
    384: T0 = 32'h9b1a06;
    385: T0 = 32'h27ffffe4;
    386: T0 = 32'hb80735d8;
    387: T0 = 32'h99be6fff;
    388: T0 = 32'h6400c5bc;
    389: T0 = 32'h26e65559;
    390: T0 = 32'h5f22d2e4;
    391: T0 = 32'hecfce58f;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T5 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T6 = reset ? 1'h0 : restartRegs_0;
  assign T7 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_14(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T5;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T6;
  reg  restartRegs_0;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (addr)
    0: T0 = 32'hcc5f16ed;
    1: T0 = 32'hb0a0f989;
    2: T0 = 32'h920d154;
    3: T0 = 32'hf7420d7;
    4: T0 = 32'hbec7e7ff;
    5: T0 = 32'ha9fffae2;
    6: T0 = 32'h42d57dbf;
    7: T0 = 32'hf0bfffa9;
    8: T0 = 32'h55cf6fff;
    9: T0 = 32'h79f4ffff;
    10: T0 = 32'hf12d757f;
    11: T0 = 32'h66b33391;
    12: T0 = 32'hd607d8;
    13: T0 = 32'hff3cc000;
    14: T0 = 32'h100f2;
    15: T0 = 32'hddf800;
    16: T0 = 32'h9100060e;
    17: T0 = 32'h17fe80;
    18: T0 = 32'h7670c3fe;
    19: T0 = 32'h20f2efc5;
    20: T0 = 32'hcbd73fff;
    21: T0 = 32'hb9fff0bb;
    22: T0 = 32'hffbe8dfe;
    23: T0 = 32'h5e3f8402;
    24: T0 = 32'hffe20f1f;
    25: T0 = 32'h5ebff440;
    26: T0 = 32'hffc0004b;
    27: T0 = 32'h113f84;
    28: T0 = 32'h9ff84606;
    29: T0 = 32'h94ff8;
    30: T0 = 32'hd97e01c8;
    31: T0 = 32'hc003f0ff;
    32: T0 = 32'hee07ea1f;
    33: T0 = 32'h700ffec7;
    34: T0 = 32'hff67bf0f;
    35: T0 = 32'ha627fffd;
    36: T0 = 32'h7ffdd6e3;
    37: T0 = 32'hab403fff;
    38: T0 = 32'h64f4cafe;
    39: T0 = 32'h5b1f7bf;
    40: T0 = 32'h11a0b81d;
    41: T0 = 32'hc010b5ff;
    42: T0 = 32'h60800205;
    43: T0 = 32'h2ec40;
    44: T0 = 32'h56024000;
    45: T0 = 32'h2400c1b4;
    46: T0 = 32'h103693c0;
    47: T0 = 32'h557cccd7;
    48: T0 = 32'hf3dbdb1;
    49: T0 = 32'h459402f;
    50: T0 = 32'hd3b8c26;
    51: T0 = 32'h828cc71f;
    52: T0 = 32'hf330727d;
    53: T0 = 32'h502bd641;
    54: T0 = 32'h3f82f119;
    55: T0 = 32'h2d745f00;
    56: T0 = 32'h5fc01b43;
    57: T0 = 32'h1fb0a80;
    58: T0 = 32'h7eec05db;
    59: T0 = 32'hc00f7198;
    60: T0 = 32'hff9101fa;
    61: T0 = 32'h5f80f78d;
    62: T0 = 32'h7ee407f;
    63: T0 = 32'h1bfefd54;
    64: T0 = 32'hf07e840f;
    65: T0 = 32'h5b9fffee;
    66: T0 = 32'hc7c37d81;
    67: T0 = 32'h17fd1ffc;
    68: T0 = 32'hf07cffef;
    69: T0 = 32'hc84361bf;
    70: T0 = 32'hbf0703fe;
    71: T0 = 32'h3ec4ffd0;
    72: T0 = 32'h39ec4007;
    73: T0 = 32'hb4f1a75;
    74: T0 = 32'h603ecf00;
    75: T0 = 32'hc2fc006f;
    76: T0 = 32'h4e61f3f8;
    77: T0 = 32'h9c018014;
    78: T0 = 32'hf62773b;
    79: T0 = 32'h14c003c0;
    80: T0 = 32'h187e0563;
    81: T0 = 32'hefa8e23e;
    82: T0 = 32'h187e07b;
    83: T0 = 32'h7cfedea1;
    84: T0 = 32'ha0380f01;
    85: T0 = 32'h87405ae0;
    86: T0 = 32'ha30301f0;
    87: T0 = 32'h10e8018c;
    88: T0 = 32'h9a08030;
    89: T0 = 32'hbe02fb;
    90: T0 = 32'hc852d41e;
    91: T0 = 32'h700fe0ed;
    92: T0 = 32'hfe8edfff;
    93: T0 = 32'h1803feef;
    94: T0 = 32'h3fe8ee4f;
    95: T0 = 32'hc6e03ffb;
    96: T0 = 32'h83ff65a8;
    97: T0 = 32'h2e9bff51;
    98: T0 = 32'heb022eef;
    99: T0 = 32'he1d50efd;
    100: T0 = 32'hf502fb2e;
    101: T0 = 32'h68ac4766;
    102: T0 = 32'h8f788a06;
    103: T0 = 32'h741001ce;
    104: T0 = 32'h29710b40;
    105: T0 = 32'hbbc18373;
    106: T0 = 32'h48b8783;
    107: T0 = 32'h57e8007f;
    108: T0 = 32'h8001f81c;
    109: T0 = 32'h55cce07;
    110: T0 = 32'hda087f91;
    111: T0 = 32'h202dc7e0;
    112: T0 = 32'hbfe207fe;
    113: T0 = 32'hc287b04f;
    114: T0 = 32'h81fff87f;
    115: T0 = 32'hfe11f96c;
    116: T0 = 32'h4876787;
    117: T0 = 32'hfbf07b2a;
    118: T0 = 32'hc0742b38;
    119: T0 = 32'hff019f;
    120: T0 = 32'hff0c2807;
    121: T0 = 32'hfb03b000;
    122: T0 = 32'h7ff01f18;
    123: T0 = 32'ha40af00;
    124: T0 = 32'h59f0147;
    125: T0 = 32'he0ea4fec;
    126: T0 = 32'h80f13800;
    127: T0 = 32'hb002a4bf;
    128: T0 = 32'h1c0f6381;
    129: T0 = 32'h7e000b48;
    130: T0 = 32'h380803c;
    131: T0 = 32'h7b8c04e;
    132: T0 = 32'h468003;
    133: T0 = 32'h603f3e02;
    134: T0 = 32'h814d5d80;
    135: T0 = 32'h830303b0;
    136: T0 = 32'h1917c74a;
    137: T0 = 32'heeb8807c;
    138: T0 = 32'h41be4e5c;
    139: T0 = 32'hfd8f7407;
    140: T0 = 32'h180ff0eb;
    141: T0 = 32'h7ff8601e;
    142: T0 = 32'ha390fd00;
    143: T0 = 32'h3fc0d99;
    144: T0 = 32'hcd221784;
    145: T0 = 32'hc1f3ba75;
    146: T0 = 32'hcf90549c;
    147: T0 = 32'h84cb80b4;
    148: T0 = 32'hf926fa1f;
    149: T0 = 32'hc41c58e0;
    150: T0 = 32'h8075f5ca;
    151: T0 = 32'h5eeed5a4;
    152: T0 = 32'h2425028b;
    153: T0 = 32'hed094bfe;
    154: T0 = 32'hac32fe15;
    155: T0 = 32'h176cdab7;
    156: T0 = 32'h53001bc6;
    157: T0 = 32'hffff0fb7;
    158: T0 = 32'hf97f7ffe;
    159: T0 = 32'he7fdc29e;
    160: T0 = 32'h8fcf01ff;
    161: T0 = 32'hc000f825;
    162: T0 = 32'h2771740f;
    163: T0 = 32'h90028602;
    164: T0 = 32'h6fd9a0;
    165: T0 = 32'he1800000;
    166: T0 = 32'h1f44a0;
    167: T0 = 32'hfe3cc0fe;
    168: T0 = 32'h3800ffea;
    169: T0 = 32'hfe8dfff;
    170: T0 = 32'h17f8ffff;
    171: T0 = 32'he1fdff5f;
    172: T0 = 32'hdb7fffbf;
    173: T0 = 32'hff1ffff7;
    174: T0 = 32'hfb0dfff9;
    175: T0 = 32'h1fbf0fed;
    176: T0 = 32'hff6e97fc;
    177: T0 = 32'hbe3803f;
    178: T0 = 32'h3fcff5f;
    179: T0 = 32'ha0fee101;
    180: T0 = 32'hf1bf0e37;
    181: T0 = 32'hfe0f9410;
    182: T0 = 32'hdf2b0032;
    183: T0 = 32'h3cfdd6c7;
    184: T0 = 32'hdff91037;
    185: T0 = 32'hdb8ef665;
    186: T0 = 32'hca8f800d;
    187: T0 = 32'h7db1015a;
    188: T0 = 32'h51331420;
    189: T0 = 32'hafe301fb;
    190: T0 = 32'h9f00;
    191: T0 = 32'h9e7eccf3;
    192: T0 = 32'hbfd1b;
    193: T0 = 32'hfc1f0133;
    194: T0 = 32'hb002d346;
    195: T0 = 32'he84eaff1;
    196: T0 = 32'he41dabeb;
    197: T0 = 32'h82a62cb2;
    198: T0 = 32'h44b79ca;
    199: T0 = 32'hacfeea6b;
    200: T0 = 32'h8c00a587;
    201: T0 = 32'h27ffbd2c;
    202: T0 = 32'hfb213710;
    203: T0 = 32'h883f036b;
    204: T0 = 32'hff83edf0;
    205: T0 = 32'h480080be;
    206: T0 = 32'h3f1fc7d;
    207: T0 = 32'ha41fc45b;
    208: T0 = 32'hf81f0359;
    209: T0 = 32'heeb13d92;
    210: T0 = 32'h7b81603b;
    211: T0 = 32'h1f758bf0;
    212: T0 = 32'hd0dc07f7;
    213: T0 = 32'he1f7fb20;
    214: T0 = 32'h7c8f003f;
    215: T0 = 32'h1e1eff40;
    216: T0 = 32'he5b08013;
    217: T0 = 32'h5df11ff8;
    218: T0 = 32'hf4f7207;
    219: T0 = 32'hd7fff8df;
    220: T0 = 32'hf07ff701;
    221: T0 = 32'he7ff1f84;
    222: T0 = 32'hfe8170cc;
    223: T0 = 32'h54107f8;
    224: T0 = 32'hec08c007;
    225: T0 = 32'h80d7c01f;
    226: T0 = 32'h2fe07e0d;
    227: T0 = 32'he2105;
    228: T0 = 32'h121e53e0;
    229: T0 = 32'h2e610748;
    230: T0 = 32'h692fee;
    231: T0 = 32'h85a6e006;
    232: T0 = 32'h70073eeb;
    233: T0 = 32'h6f88ff02;
    234: T0 = 32'h682504bf;
    235: T0 = 32'hc730fdc8;
    236: T0 = 32'h3c02e;
    237: T0 = 32'h1ea4a7f4;
    238: T0 = 32'hb0000a0c;
    239: T0 = 32'hbecd78bd;
    240: T0 = 32'hce007f90;
    241: T0 = 32'h37349f13;
    242: T0 = 32'h8d03bfd;
    243: T0 = 32'h5600a0ae;
    244: T0 = 32'h10412aa3;
    245: T0 = 32'h6023754b;
    246: T0 = 32'h30ec3e21;
    247: T0 = 32'hce551256;
    248: T0 = 32'h8a6ab9cb;
    249: T0 = 32'h627b42d9;
    250: T0 = 32'h8881eab8;
    251: T0 = 32'h1cf279f;
    252: T0 = 32'h6c801db4;
    253: T0 = 32'h400e1c4;
    254: T0 = 32'he0c07fe2;
    255: T0 = 32'hff1e7aff;
    256: T0 = 32'hf64afff8;
    257: T0 = 32'h300cd3;
    258: T0 = 32'h5400f8e;
    259: T0 = 32'hc03e;
    260: T0 = 32'h40d800;
    261: T0 = 32'he4001801;
    262: T0 = 32'hf01a0ac0;
    263: T0 = 32'hb81d03c0;
    264: T0 = 32'hffff0119;
    265: T0 = 32'hff7b38fc;
    266: T0 = 32'hdfffc47e;
    267: T0 = 32'hfff15c0f;
    268: T0 = 32'ha9ffe623;
    269: T0 = 32'he1ff1a01;
    270: T0 = 32'hf9bf1040;
    271: T0 = 32'hf00b0150;
    272: T0 = 32'h96b8c000;
    273: T0 = 32'h86142025;
    274: T0 = 32'h1f257c08;
    275: T0 = 32'h60200603;
    276: T0 = 32'h3e03f80;
    277: T0 = 32'h27c410f0;
    278: T0 = 32'h403efd4b;
    279: T0 = 32'hea649e9f;
    280: T0 = 32'h1003fffa;
    281: T0 = 32'hf481f7ff;
    282: T0 = 32'h247fdff;
    283: T0 = 32'hfc0ff23f;
    284: T0 = 32'hc77dff8f;
    285: T0 = 32'h7fee5e27;
    286: T0 = 32'h3c0e67fb;
    287: T0 = 32'hf7ff4009;
    288: T0 = 32'h91b2b286;
    289: T0 = 32'hcf5f8000;
    290: T0 = 32'hec0c1ccd;
    291: T0 = 32'hdec3b061;
    292: T0 = 32'he8833a6a;
    293: T0 = 32'hdcc1f70b;
    294: T0 = 32'h7edf9bc4;
    295: T0 = 32'hc482f79b;
    296: T0 = 32'hf4e3d6d6;
    297: T0 = 32'hcf48754e;
    298: T0 = 32'h271020a;
    299: T0 = 32'h5ffaef46;
    300: T0 = 32'ha17d0107;
    301: T0 = 32'h26f93eec;
    302: T0 = 32'h6478810;
    303: T0 = 32'h11680408;
    304: T0 = 32'hffc0bb40;
    305: T0 = 32'h187f00b4;
    306: T0 = 32'h7fff02a1;
    307: T0 = 32'he07d600e;
    308: T0 = 32'h8bff037d;
    309: T0 = 32'h566f70;
    310: T0 = 32'hb000fc13;
    311: T0 = 32'h2603ff;
    312: T0 = 32'h4f00ffe0;
    313: T0 = 32'h18877;
    314: T0 = 32'h1010ffff;
    315: T0 = 32'h8e00fe9b;
    316: T0 = 32'h95f2fb;
    317: T0 = 32'h53fc5fe1;
    318: T0 = 32'hcff9f53f;
    319: T0 = 32'hd01fefff;
    320: T0 = 32'hf0fffec7;
    321: T0 = 32'hfe167fff;
    322: T0 = 32'hf41ffff5;
    323: T0 = 32'hffc380df;
    324: T0 = 32'h6d83ffff;
    325: T0 = 32'h1ff8fe46;
    326: T0 = 32'hda0bfff;
    327: T0 = 32'h8f76f89d;
    328: T0 = 32'hdfe01f;
    329: T0 = 32'h39780484;
    330: T0 = 32'h8013100c;
    331: T0 = 32'hd38c0000;
    332: T0 = 32'hff47e042;
    333: T0 = 32'hfacc0080;
    334: T0 = 32'ha90f049d;
    335: T0 = 32'hff1e6b8f;
    336: T0 = 32'hdf970276;
    337: T0 = 32'h3ffa3e00;
    338: T0 = 32'hf4fc0186;
    339: T0 = 32'hc0021378;
    340: T0 = 32'h5e43010;
    341: T0 = 32'hdae84ce9;
    342: T0 = 32'h7a4dccd8;
    343: T0 = 32'h1ce6c8b2;
    344: T0 = 32'h5acf408a;
    345: T0 = 32'h49764aea;
    346: T0 = 32'h2dc3978e;
    347: T0 = 32'h7ab89c0f;
    348: T0 = 32'h7cd70297;
    349: T0 = 32'hf1bc100;
    350: T0 = 32'hbffc8012;
    351: T0 = 32'h4077e749;
    352: T0 = 32'hcff0001;
    353: T0 = 32'h80177f60;
    354: T0 = 32'he30f0f80;
    355: T0 = 32'h68000f8c;
    356: T0 = 32'h3f444bfc;
    357: T0 = 32'h70f025;
    358: T0 = 32'h83f505df;
    359: T0 = 32'h8803ffe3;
    360: T0 = 32'h753833f;
    361: T0 = 32'hba00ffff;
    362: T0 = 32'h2bcfc27;
    363: T0 = 32'hf3d8ff86;
    364: T0 = 32'h81fb07e3;
    365: T0 = 32'h1f1b4be0;
    366: T0 = 32'hd03f0425;
    367: T0 = 32'hf1f037ee;
    368: T0 = 32'h8403a064;
    369: T0 = 32'h3f0dc96d;
    370: T0 = 32'hf874b801;
    371: T0 = 32'hc3f80f64;
    372: T0 = 32'h8f0b2a00;
    373: T0 = 32'hdc1f20fc;
    374: T0 = 32'hfcf0a618;
    375: T0 = 32'h100c00f;
    376: T0 = 32'h7fcfd12;
    377: T0 = 32'h81646201;
    378: T0 = 32'ha0001fe1;
    379: T0 = 32'h701d4800;
    380: T0 = 32'h2400c3c6;
    381: T0 = 32'h1f83f682;
    382: T0 = 32'h3ac67f8;
    383: T0 = 32'h80dfe8;
    384: T0 = 32'h7cccc0af;
    385: T0 = 32'h240e0b1;
    386: T0 = 32'h283c587;
    387: T0 = 32'h5d4b7fbc;
    388: T0 = 32'h1fd05d4c;
    389: T0 = 32'he4885fff;
    390: T0 = 32'hc087af99;
    391: T0 = 32'hf2620edd;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T5 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T6 = reset ? 1'h0 : restartRegs_0;
  assign T7 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_15(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T5;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T6;
  reg  restartRegs_0;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (addr)
    0: T0 = 32'hf37a9bc8;
    1: T0 = 32'h334d44a3;
    2: T0 = 32'hd75be605;
    3: T0 = 32'h14f1714e;
    4: T0 = 32'hf56ca004;
    5: T0 = 32'h228c2ed0;
    6: T0 = 32'hf982a6f3;
    7: T0 = 32'h16038155;
    8: T0 = 32'h7ff7ae7f;
    9: T0 = 32'hadc0f831;
    10: T0 = 32'h1ffd535b;
    11: T0 = 32'h61b03f00;
    12: T0 = 32'hc1f86dd9;
    13: T0 = 32'hd098f0;
    14: T0 = 32'hd81f025e;
    15: T0 = 32'he0093b8f;
    16: T0 = 32'hffc1781c;
    17: T0 = 32'he002438;
    18: T0 = 32'h5883f8;
    19: T0 = 32'he0f0c14f;
    20: T0 = 32'hfec9981f;
    21: T0 = 32'hbd0fff83;
    22: T0 = 32'hfff13c00;
    23: T0 = 32'hfd4803fd;
    24: T0 = 32'h8fff73e0;
    25: T0 = 32'hf4fe401f;
    26: T0 = 32'he47fffe5;
    27: T0 = 32'h3e17fa00;
    28: T0 = 32'h7f150380;
    29: T0 = 32'h7ff03bf4;
    30: T0 = 32'hcbfdc03e;
    31: T0 = 32'hf7fce09f;
    32: T0 = 32'h3ff3907;
    33: T0 = 32'hb0477275;
    34: T0 = 32'hc02687e0;
    35: T0 = 32'h10818f25;
    36: T0 = 32'hb08260fe;
    37: T0 = 32'hc40c68f4;
    38: T0 = 32'h57ab0ea5;
    39: T0 = 32'h14616db8;
    40: T0 = 32'h817edc04;
    41: T0 = 32'hd03257d6;
    42: T0 = 32'h482f9bab;
    43: T0 = 32'hef4480ed;
    44: T0 = 32'h82ff486e;
    45: T0 = 32'hf00d0b30;
    46: T0 = 32'hd3670100;
    47: T0 = 32'h3e82f94c;
    48: T0 = 32'hcbba2391;
    49: T0 = 32'had281779;
    50: T0 = 32'h2b9cc5f;
    51: T0 = 32'h77ab7668;
    52: T0 = 32'h4495c6a0;
    53: T0 = 32'h66017be4;
    54: T0 = 32'hd4461af8;
    55: T0 = 32'h6d25213e;
    56: T0 = 32'hcd8060de;
    57: T0 = 32'h3e0f9742;
    58: T0 = 32'hd80fdd2;
    59: T0 = 32'hff9582f;
    60: T0 = 32'haf107ff0;
    61: T0 = 32'h3ff04f0;
    62: T0 = 32'hf7daa03e;
    63: T0 = 32'h607f00ac;
    64: T0 = 32'hfff1fa00;
    65: T0 = 32'h860f0008;
    66: T0 = 32'hffc7b701;
    67: T0 = 32'h3dc1fc19;
    68: T0 = 32'h1ff8fbb0;
    69: T0 = 32'h66bfff;
    70: T0 = 32'he1f8fff2;
    71: T0 = 32'h41fff;
    72: T0 = 32'h660ffffe;
    73: T0 = 32'hf000f1ff;
    74: T0 = 32'h4e0ffff;
    75: T0 = 32'h700ff87;
    76: T0 = 32'h4047df79;
    77: T0 = 32'h783987ff;
    78: T0 = 32'h1f80b5bf;
    79: T0 = 32'h65f3f01f;
    80: T0 = 32'h33f8fabf;
    81: T0 = 32'hcdcffe00;
    82: T0 = 32'h5d0f43f3;
    83: T0 = 32'h7c85adc0;
    84: T0 = 32'hbe440411;
    85: T0 = 32'h4386bfbc;
    86: T0 = 32'he48200e6;
    87: T0 = 32'hd8180a3b;
    88: T0 = 32'h83b00036;
    89: T0 = 32'h741d84eb;
    90: T0 = 32'h210b0463;
    91: T0 = 32'h8fbf9017;
    92: T0 = 32'h2c239107;
    93: T0 = 32'h5644ca04;
    94: T0 = 32'hffe71ac5;
    95: T0 = 32'hd625c833;
    96: T0 = 32'hb65f474c;
    97: T0 = 32'h1fade0bb;
    98: T0 = 32'hf36d8aac;
    99: T0 = 32'h81ef9585;
    100: T0 = 32'h678a6c38;
    101: T0 = 32'hc8c93e8;
    102: T0 = 32'hb9f5726b;
    103: T0 = 32'hd4a94eeb;
    104: T0 = 32'hd034f601;
    105: T0 = 32'h97f825bc;
    106: T0 = 32'h90069f8;
    107: T0 = 32'h8ea8fffa;
    108: T0 = 32'h7f953f;
    109: T0 = 32'hf938fe3f;
    110: T0 = 32'h8007bac3;
    111: T0 = 32'h1fe99fc0;
    112: T0 = 32'he80002a7;
    113: T0 = 32'hc07837ff;
    114: T0 = 32'h889ff05f;
    115: T0 = 32'hfe0761bf;
    116: T0 = 32'h2de78f02;
    117: T0 = 32'h1fe01187;
    118: T0 = 32'h3407838;
    119: T0 = 32'hc0ff3e19;
    120: T0 = 32'hfc1f6b01;
    121: T0 = 32'hba0703d0;
    122: T0 = 32'hf3f9d478;
    123: T0 = 32'hb243017e;
    124: T0 = 32'h3f9febed;
    125: T0 = 32'hc14cf043;
    126: T0 = 32'h87f93a75;
    127: T0 = 32'h35360c;
    128: T0 = 32'h823f21ff;
    129: T0 = 32'hf803e570;
    130: T0 = 32'h7e44df0f;
    131: T0 = 32'h2780fe8f;
    132: T0 = 32'h78cec50;
    133: T0 = 32'h15c0fec;
    134: T0 = 32'he0f770fd;
    135: T0 = 32'h7207e8fe;
    136: T0 = 32'hc3e7e63f;
    137: T0 = 32'h5820ffff;
    138: T0 = 32'h1621fe56;
    139: T0 = 32'hf1838fff;
    140: T0 = 32'h58c0fa35;
    141: T0 = 32'h4fa20349;
    142: T0 = 32'h43520001;
    143: T0 = 32'hedeb9344;
    144: T0 = 32'h7fa40000;
    145: T0 = 32'h47ea3362;
    146: T0 = 32'h22a17981;
    147: T0 = 32'h486f37cc;
    148: T0 = 32'hc0891f7e;
    149: T0 = 32'he717a5b;
    150: T0 = 32'hbaf32f64;
    151: T0 = 32'h41dea804;
    152: T0 = 32'h8406e332;
    153: T0 = 32'he41c7d01;
    154: T0 = 32'hb0111f9b;
    155: T0 = 32'h77fe09c0;
    156: T0 = 32'h47000ffb;
    157: T0 = 32'hdbf2a78;
    158: T0 = 32'hd4f883f8;
    159: T0 = 32'hc02fcb85;
    160: T0 = 32'hbe6fc03f;
    161: T0 = 32'hbf01fd20;
    162: T0 = 32'he1f6d80f;
    163: T0 = 32'he3ffffff;
    164: T0 = 32'hfe0ff5a1;
    165: T0 = 32'hfc3f1f7f;
    166: T0 = 32'hffe0ff0a;
    167: T0 = 32'h7c741f0;
    168: T0 = 32'hbcbc81f9;
    169: T0 = 32'hc07cf00f;
    170: T0 = 32'hbbc10c07;
    171: T0 = 32'h340f2d00;
    172: T0 = 32'hfabc0380;
    173: T0 = 32'hcc4000cf;
    174: T0 = 32'h1fbf7870;
    175: T0 = 32'hbca81c07;
    176: T0 = 32'hc3f647b7;
    177: T0 = 32'hcfca21e0;
    178: T0 = 32'hfc3f0a5e;
    179: T0 = 32'hecfce49f;
    180: T0 = 32'hc8e3f026;
    181: T0 = 32'hecfbe8c;
    182: T0 = 32'h1dce4703;
    183: T0 = 32'h41fd2fd9;
    184: T0 = 32'h93dc0c60;
    185: T0 = 32'h753f01ea;
    186: T0 = 32'he1dfe078;
    187: T0 = 32'hff07817d;
    188: T0 = 32'hfd0a1fd3;
    189: T0 = 32'h2f809803;
    190: T0 = 32'h4b07f3b7;
    191: T0 = 32'h9f8ff80;
    192: T0 = 32'h80001090;
    193: T0 = 32'h3a0bdffc;
    194: T0 = 32'hb8002d5a;
    195: T0 = 32'hfe5b677d;
    196: T0 = 32'h91b5c930;
    197: T0 = 32'hca940f22;
    198: T0 = 32'hd5a64930;
    199: T0 = 32'hab95877a;
    200: T0 = 32'h5ec2d66;
    201: T0 = 32'h143fb9b;
    202: T0 = 32'h37186bb;
    203: T0 = 32'hf0005fe3;
    204: T0 = 32'hbfce10c0;
    205: T0 = 32'h5f0c18ff;
    206: T0 = 32'hdfe5ee7c;
    207: T0 = 32'h7f0c3e1;
    208: T0 = 32'h8400032f;
    209: T0 = 32'hb7881f;
    210: T0 = 32'h9780e41d;
    211: T0 = 32'h80832f01;
    212: T0 = 32'hb7ff0f13;
    213: T0 = 32'hffce1278;
    214: T0 = 32'hf19f007e;
    215: T0 = 32'hfffffb78;
    216: T0 = 32'hfe774003;
    217: T0 = 32'h7fef1fe0;
    218: T0 = 32'h3ff72010;
    219: T0 = 32'h340ec0ff;
    220: T0 = 32'h40fef468;
    221: T0 = 32'h2886a007;
    222: T0 = 32'h20003fde;
    223: T0 = 32'h37bfe0;
    224: T0 = 32'h770007f3;
    225: T0 = 32'h1eabfe;
    226: T0 = 32'hcc38fc07;
    227: T0 = 32'ha002367f;
    228: T0 = 32'h7c007fc0;
    229: T0 = 32'h63010a11;
    230: T0 = 32'hff49b7ce;
    231: T0 = 32'hc08ff0a2;
    232: T0 = 32'h7ff98b6d;
    233: T0 = 32'h80b9705;
    234: T0 = 32'h4ffd079b;
    235: T0 = 32'hbe4020dc;
    236: T0 = 32'h27f6e039;
    237: T0 = 32'h27f339;
    238: T0 = 32'hb078cf0b;
    239: T0 = 32'h142e;
    240: T0 = 32'hf4bbe1f0;
    241: T0 = 32'hfc02d7a5;
    242: T0 = 32'h1006afb6;
    243: T0 = 32'h27b217fe;
    244: T0 = 32'h94e1fe0e;
    245: T0 = 32'h45546f7;
    246: T0 = 32'h95640e3a;
    247: T0 = 32'h54911abc;
    248: T0 = 32'ha63334e6;
    249: T0 = 32'h1a1ecb49;
    250: T0 = 32'hfe7b7c0f;
    251: T0 = 32'h9b631259;
    252: T0 = 32'h71851ee2;
    253: T0 = 32'he367bf67;
    254: T0 = 32'h10005af6;
    255: T0 = 32'hc27f730;
    256: T0 = 32'h4f30db2d;
    257: T0 = 32'h818bb743;
    258: T0 = 32'hb31a7ff;
    259: T0 = 32'h7e009747;
    260: T0 = 32'he2df6401;
    261: T0 = 32'h5bff01ea;
    262: T0 = 32'hfe07c2c0;
    263: T0 = 32'h123f001f;
    264: T0 = 32'hfff0d80c;
    265: T0 = 32'ha3c03f;
    266: T0 = 32'h7f8fffc2;
    267: T0 = 32'hf805fe3f;
    268: T0 = 32'h9b21fff8;
    269: T0 = 32'h3fc00715;
    270: T0 = 32'hd9097fe;
    271: T0 = 32'h1fc80fd;
    272: T0 = 32'h4aaadf;
    273: T0 = 32'h531f000c;
    274: T0 = 32'he2174180;
    275: T0 = 32'hb2990000;
    276: T0 = 32'h1f72397a;
    277: T0 = 32'hf7d08100;
    278: T0 = 32'he0f80f8b;
    279: T0 = 32'hfa86ba08;
    280: T0 = 32'hcf8f47fe;
    281: T0 = 32'h7de62e82;
    282: T0 = 32'habc0bff;
    283: T0 = 32'h87ede942;
    284: T0 = 32'hd72c00ff;
    285: T0 = 32'h243fa0ac;
    286: T0 = 32'hfd0f9003;
    287: T0 = 32'h42020c81;
    288: T0 = 32'hcf8c8002;
    289: T0 = 32'h8a002655;
    290: T0 = 32'he7dbf04;
    291: T0 = 32'h40600f5f;
    292: T0 = 32'ha4713669;
    293: T0 = 32'h206727b2;
    294: T0 = 32'h81ac1305;
    295: T0 = 32'hb4008e06;
    296: T0 = 32'h611b7e8d;
    297: T0 = 32'hfd27f7ca;
    298: T0 = 32'h3c9ae190;
    299: T0 = 32'hf90103ad;
    300: T0 = 32'h1aeed950;
    301: T0 = 32'h3e80c00f;
    302: T0 = 32'h3fa3b9f;
    303: T0 = 32'h1ff0ff80;
    304: T0 = 32'h56364b;
    305: T0 = 32'hfdf8fffc;
    306: T0 = 32'hfc07518f;
    307: T0 = 32'h27ebfe5d;
    308: T0 = 32'h7fe0d37d;
    309: T0 = 32'h80f36bff;
    310: T0 = 32'hdfff7c4f;
    311: T0 = 32'hfe02183f;
    312: T0 = 32'hdafe0c0;
    313: T0 = 32'hfbf004ff;
    314: T0 = 32'h60fc06;
    315: T0 = 32'hf720c;
    316: T0 = 32'hfc020b80;
    317: T0 = 32'h241807ea;
    318: T0 = 32'he7204780;
    319: T0 = 32'h94600078;
    320: T0 = 32'he7ed114;
    321: T0 = 32'hffa0c003;
    322: T0 = 32'h41f73a3b;
    323: T0 = 32'hc7fa6480;
    324: T0 = 32'ha44f0027;
    325: T0 = 32'h7c3de95c;
    326: T0 = 32'hc719fc16;
    327: T0 = 32'h31c3ffaf;
    328: T0 = 32'h1e0c3fe1;
    329: T0 = 32'h800ebffb;
    330: T0 = 32'h41e2f3ff;
    331: T0 = 32'hb90cfffe;
    332: T0 = 32'ha39ff82f;
    333: T0 = 32'hff02ffff;
    334: T0 = 32'h199fe7ff;
    335: T0 = 32'h7d07efff;
    336: T0 = 32'ha020fa14;
    337: T0 = 32'h8f4edf23;
    338: T0 = 32'h3c00fa00;
    339: T0 = 32'h1e2b29e;
    340: T0 = 32'h64c07f52;
    341: T0 = 32'h901e3281;
    342: T0 = 32'h6ad60b72;
    343: T0 = 32'h8b2126fd;
    344: T0 = 32'hfa57eb7b;
    345: T0 = 32'hc2fef76e;
    346: T0 = 32'h874607f0;
    347: T0 = 32'hb0f4be35;
    348: T0 = 32'hc4ff59b1;
    349: T0 = 32'hf2d09480;
    350: T0 = 32'h1bf03af;
    351: T0 = 32'hffed1460;
    352: T0 = 32'h17bf3982;
    353: T0 = 32'h1fffc44c;
    354: T0 = 32'hc55e003f;
    355: T0 = 32'hf15f7f98;
    356: T0 = 32'hff6b4800;
    357: T0 = 32'hffff0222;
    358: T0 = 32'hfdf7abe0;
    359: T0 = 32'heb7f7007;
    360: T0 = 32'hff00389f;
    361: T0 = 32'h1691f3fe;
    362: T0 = 32'h380ffa7;
    363: T0 = 32'h78189f;
    364: T0 = 32'h80603ff1;
    365: T0 = 32'h1e4c09;
    366: T0 = 32'he00e01ff;
    367: T0 = 32'h6000fe87;
    368: T0 = 32'h1f005e3f;
    369: T0 = 32'hd02af24;
    370: T0 = 32'hdc43ff;
    371: T0 = 32'hc8f00d;
    372: T0 = 32'h55827;
    373: T0 = 32'h3a162e00;
    374: T0 = 32'h200007a0;
    375: T0 = 32'h3ee00000;
    376: T0 = 32'ha180003b;
    377: T0 = 32'hf0a7900;
    378: T0 = 32'h27fe000f;
    379: T0 = 32'hfff97cde;
    380: T0 = 32'he5ff5021;
    381: T0 = 32'hfffffaf7;
    382: T0 = 32'hf9bff37f;
    383: T0 = 32'hde1fffab;
    384: T0 = 32'h89db5103;
    385: T0 = 32'h5f0867e2;
    386: T0 = 32'hfdf567b1;
    387: T0 = 32'h6905144a;
    388: T0 = 32'hbfff7008;
    389: T0 = 32'h70c30000;
    390: T0 = 32'h9fffcac3;
    391: T0 = 32'hfa82f57;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T5 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T6 = reset ? 1'h0 : restartRegs_0;
  assign T7 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_16(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[7:0] io_weights
);

  reg [7:0] weightsReg;
  wire[7:0] T4;
  reg [7:0] T0;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T5;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T6;
  reg  restartRegs_0;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 8'h0 : T0;
  always @(*) case (addr)
    0: T0 = 8'hd;
    1: T0 = 8'h1a;
    2: T0 = 8'h14;
    3: T0 = 8'h18;
    4: T0 = 8'he3;
    5: T0 = 8'he8;
    6: T0 = 8'hc9;
    7: T0 = 8'h39;
    8: T0 = 8'hce;
    9: T0 = 8'hee;
    10: T0 = 8'hd3;
    11: T0 = 8'h18;
    12: T0 = 8'h0;
    13: T0 = 8'hd7;
    14: T0 = 8'h6;
    15: T0 = 8'hf9;
    16: T0 = 8'h0;
    17: T0 = 8'h23;
    18: T0 = 8'heb;
    19: T0 = 8'h11;
    20: T0 = 8'he9;
    21: T0 = 8'h2a;
    22: T0 = 8'h1;
    23: T0 = 8'hfd;
    24: T0 = 8'hd;
    25: T0 = 8'hde;
    26: T0 = 8'hfd;
    27: T0 = 8'hcc;
    28: T0 = 8'h33;
    29: T0 = 8'he4;
    30: T0 = 8'hf3;
    31: T0 = 8'hf;
    32: T0 = 8'h0;
    33: T0 = 8'h0;
    34: T0 = 8'h0;
    35: T0 = 8'h0;
    36: T0 = 8'h0;
    37: T0 = 8'h0;
    38: T0 = 8'h0;
    39: T0 = 8'h0;
    40: T0 = 8'h0;
    41: T0 = 8'h0;
    42: T0 = 8'h0;
    43: T0 = 8'h0;
    44: T0 = 8'h0;
    45: T0 = 8'h0;
    46: T0 = 8'h0;
    47: T0 = 8'h0;
    48: T0 = 8'h0;
    49: T0 = 8'h6;
    50: T0 = 8'hd4;
    51: T0 = 8'hc6;
    52: T0 = 8'hdd;
    53: T0 = 8'hf6;
    54: T0 = 8'hdc;
    55: T0 = 8'hb;
    56: T0 = 8'h8;
    57: T0 = 8'he8;
    58: T0 = 8'hdf;
    59: T0 = 8'h9;
    60: T0 = 8'hdc;
    61: T0 = 8'h8;
    62: T0 = 8'he7;
    63: T0 = 8'hef;
    64: T0 = 8'h23;
    65: T0 = 8'hd8;
    66: T0 = 8'hf7;
    67: T0 = 8'he3;
    68: T0 = 8'h3f;
    69: T0 = 8'h6;
    70: T0 = 8'hf4;
    71: T0 = 8'hf8;
    72: T0 = 8'h3;
    73: T0 = 8'he1;
    74: T0 = 8'h3d;
    75: T0 = 8'hf0;
    76: T0 = 8'h20;
    77: T0 = 8'h7;
    78: T0 = 8'hec;
    79: T0 = 8'h1a;
    80: T0 = 8'hef;
    81: T0 = 8'h0;
    82: T0 = 8'h0;
    83: T0 = 8'h0;
    84: T0 = 8'h0;
    85: T0 = 8'h0;
    86: T0 = 8'h0;
    87: T0 = 8'h0;
    88: T0 = 8'h0;
    89: T0 = 8'h0;
    90: T0 = 8'h0;
    91: T0 = 8'h0;
    92: T0 = 8'h0;
    93: T0 = 8'h0;
    94: T0 = 8'h0;
    95: T0 = 8'h0;
    96: T0 = 8'h0;
    97: T0 = 8'h0;
    98: T0 = 8'heb;
    99: T0 = 8'hd9;
    100: T0 = 8'h1e;
    101: T0 = 8'hfd;
    102: T0 = 8'h36;
    103: T0 = 8'h27;
    104: T0 = 8'hfd;
    105: T0 = 8'hf1;
    106: T0 = 8'he7;
    107: T0 = 8'h19;
    108: T0 = 8'h9;
    109: T0 = 8'h1;
    110: T0 = 8'h8;
    111: T0 = 8'hf2;
    112: T0 = 8'h3f;
    113: T0 = 8'hf1;
    114: T0 = 8'hf9;
    115: T0 = 8'hd7;
    116: T0 = 8'hf9;
    117: T0 = 8'hd0;
    118: T0 = 8'hf4;
    119: T0 = 8'hc9;
    120: T0 = 8'hb;
    121: T0 = 8'h10;
    122: T0 = 8'hfa;
    123: T0 = 8'h3f;
    124: T0 = 8'hec;
    125: T0 = 8'h30;
    126: T0 = 8'hdc;
    127: T0 = 8'hd3;
    128: T0 = 8'h1a;
    129: T0 = 8'hea;
    130: T0 = 8'h0;
    131: T0 = 8'h0;
    132: T0 = 8'h0;
    133: T0 = 8'h0;
    134: T0 = 8'h0;
    135: T0 = 8'h0;
    136: T0 = 8'h0;
    137: T0 = 8'h0;
    138: T0 = 8'h0;
    139: T0 = 8'h0;
    140: T0 = 8'h0;
    141: T0 = 8'h0;
    142: T0 = 8'h0;
    143: T0 = 8'h0;
    144: T0 = 8'h0;
    145: T0 = 8'h0;
    146: T0 = 8'h0;
    147: T0 = 8'hea;
    148: T0 = 8'h21;
    149: T0 = 8'ha;
    150: T0 = 8'h6;
    151: T0 = 8'hea;
    152: T0 = 8'hed;
    153: T0 = 8'hef;
    154: T0 = 8'hf0;
    155: T0 = 8'hb;
    156: T0 = 8'h9;
    157: T0 = 8'hd;
    158: T0 = 8'ha;
    159: T0 = 8'he;
    160: T0 = 8'h8;
    161: T0 = 8'h22;
    162: T0 = 8'h2;
    163: T0 = 8'he0;
    164: T0 = 8'hc0;
    165: T0 = 8'hfb;
    166: T0 = 8'hff;
    167: T0 = 8'heb;
    168: T0 = 8'hfa;
    169: T0 = 8'hdd;
    170: T0 = 8'h1f;
    171: T0 = 8'h23;
    172: T0 = 8'hfa;
    173: T0 = 8'he9;
    174: T0 = 8'hff;
    175: T0 = 8'h21;
    176: T0 = 8'h19;
    177: T0 = 8'hf1;
    178: T0 = 8'h2c;
    179: T0 = 8'h0;
    180: T0 = 8'h0;
    181: T0 = 8'h0;
    182: T0 = 8'h0;
    183: T0 = 8'h0;
    184: T0 = 8'h0;
    185: T0 = 8'h0;
    186: T0 = 8'h0;
    187: T0 = 8'h0;
    188: T0 = 8'h0;
    189: T0 = 8'h0;
    190: T0 = 8'h0;
    191: T0 = 8'h0;
    192: T0 = 8'h0;
    193: T0 = 8'h0;
    194: T0 = 8'h0;
    195: T0 = 8'h0;
    196: T0 = 8'hd7;
    197: T0 = 8'h5;
    198: T0 = 8'hf2;
    199: T0 = 8'h6;
    200: T0 = 8'hf7;
    201: T0 = 8'h27;
    202: T0 = 8'hf8;
    203: T0 = 8'hcf;
    204: T0 = 8'h25;
    205: T0 = 8'h1b;
    206: T0 = 8'hfe;
    207: T0 = 8'h13;
    208: T0 = 8'hec;
    209: T0 = 8'he5;
    210: T0 = 8'hd;
    211: T0 = 8'h2b;
    212: T0 = 8'h3;
    213: T0 = 8'hd;
    214: T0 = 8'hd6;
    215: T0 = 8'hf1;
    216: T0 = 8'hd2;
    217: T0 = 8'hf1;
    218: T0 = 8'h12;
    219: T0 = 8'h18;
    220: T0 = 8'h11;
    221: T0 = 8'hd4;
    222: T0 = 8'he1;
    223: T0 = 8'h4;
    224: T0 = 8'h4;
    225: T0 = 8'he6;
    226: T0 = 8'hc;
    227: T0 = 8'he2;
    228: T0 = 8'h0;
    229: T0 = 8'h0;
    230: T0 = 8'h0;
    231: T0 = 8'h0;
    232: T0 = 8'h0;
    233: T0 = 8'h0;
    234: T0 = 8'h0;
    235: T0 = 8'h0;
    236: T0 = 8'h0;
    237: T0 = 8'h0;
    238: T0 = 8'h0;
    239: T0 = 8'h0;
    240: T0 = 8'h0;
    241: T0 = 8'h0;
    242: T0 = 8'h0;
    243: T0 = 8'h0;
    244: T0 = 8'h0;
    245: T0 = 8'he;
    246: T0 = 8'h17;
    247: T0 = 8'hb;
    248: T0 = 8'h22;
    249: T0 = 8'hf8;
    250: T0 = 8'h5;
    251: T0 = 8'hf8;
    252: T0 = 8'hee;
    253: T0 = 8'hec;
    254: T0 = 8'h16;
    255: T0 = 8'he4;
    256: T0 = 8'h19;
    257: T0 = 8'h19;
    258: T0 = 8'h4;
    259: T0 = 8'h8;
    260: T0 = 8'he7;
    261: T0 = 8'hfd;
    262: T0 = 8'h1;
    263: T0 = 8'hef;
    264: T0 = 8'hee;
    265: T0 = 8'hed;
    266: T0 = 8'hee;
    267: T0 = 8'hce;
    268: T0 = 8'h17;
    269: T0 = 8'hcf;
    270: T0 = 8'h17;
    271: T0 = 8'hd7;
    272: T0 = 8'h39;
    273: T0 = 8'hec;
    274: T0 = 8'h3;
    275: T0 = 8'he2;
    276: T0 = 8'hfb;
    277: T0 = 8'h0;
    278: T0 = 8'h0;
    279: T0 = 8'h0;
    280: T0 = 8'h0;
    281: T0 = 8'h0;
    282: T0 = 8'h0;
    283: T0 = 8'h0;
    284: T0 = 8'h0;
    285: T0 = 8'h0;
    286: T0 = 8'h0;
    287: T0 = 8'h0;
    288: T0 = 8'h0;
    289: T0 = 8'h0;
    290: T0 = 8'h0;
    291: T0 = 8'h0;
    292: T0 = 8'h0;
    293: T0 = 8'h0;
    294: T0 = 8'h24;
    295: T0 = 8'h13;
    296: T0 = 8'h0;
    297: T0 = 8'h4;
    298: T0 = 8'h36;
    299: T0 = 8'he1;
    300: T0 = 8'hfc;
    301: T0 = 8'h13;
    302: T0 = 8'h3f;
    303: T0 = 8'hf;
    304: T0 = 8'h21;
    305: T0 = 8'h2c;
    306: T0 = 8'h16;
    307: T0 = 8'h5;
    308: T0 = 8'h32;
    309: T0 = 8'h11;
    310: T0 = 8'h2b;
    311: T0 = 8'h28;
    312: T0 = 8'hd;
    313: T0 = 8'hc0;
    314: T0 = 8'hd5;
    315: T0 = 8'h24;
    316: T0 = 8'hb;
    317: T0 = 8'hc0;
    318: T0 = 8'hdb;
    319: T0 = 8'hfc;
    320: T0 = 8'h27;
    321: T0 = 8'hfe;
    322: T0 = 8'h2;
    323: T0 = 8'hb;
    324: T0 = 8'h26;
    325: T0 = 8'hf1;
    326: T0 = 8'h0;
    327: T0 = 8'h0;
    328: T0 = 8'h0;
    329: T0 = 8'h0;
    330: T0 = 8'h0;
    331: T0 = 8'h0;
    332: T0 = 8'h0;
    333: T0 = 8'h0;
    334: T0 = 8'h0;
    335: T0 = 8'h0;
    336: T0 = 8'h0;
    337: T0 = 8'h0;
    338: T0 = 8'h0;
    339: T0 = 8'h0;
    340: T0 = 8'h0;
    341: T0 = 8'h0;
    342: T0 = 8'h0;
    343: T0 = 8'hc;
    344: T0 = 8'hd2;
    345: T0 = 8'h14;
    346: T0 = 8'hfa;
    347: T0 = 8'hdb;
    348: T0 = 8'hf9;
    349: T0 = 8'hf;
    350: T0 = 8'hf4;
    351: T0 = 8'hff;
    352: T0 = 8'h1b;
    353: T0 = 8'hfc;
    354: T0 = 8'h1;
    355: T0 = 8'hfa;
    356: T0 = 8'h8;
    357: T0 = 8'hda;
    358: T0 = 8'h6;
    359: T0 = 8'h4;
    360: T0 = 8'h28;
    361: T0 = 8'hfc;
    362: T0 = 8'h0;
    363: T0 = 8'h33;
    364: T0 = 8'hed;
    365: T0 = 8'h3f;
    366: T0 = 8'hd1;
    367: T0 = 8'hfb;
    368: T0 = 8'hf8;
    369: T0 = 8'h14;
    370: T0 = 8'h3f;
    371: T0 = 8'hf4;
    372: T0 = 8'hd5;
    373: T0 = 8'hef;
    374: T0 = 8'h19;
    375: T0 = 8'h0;
    376: T0 = 8'h0;
    377: T0 = 8'h0;
    378: T0 = 8'h0;
    379: T0 = 8'h0;
    380: T0 = 8'h0;
    381: T0 = 8'h0;
    382: T0 = 8'h0;
    383: T0 = 8'h0;
    384: T0 = 8'h0;
    385: T0 = 8'h0;
    386: T0 = 8'h0;
    387: T0 = 8'h0;
    388: T0 = 8'h0;
    389: T0 = 8'h0;
    390: T0 = 8'h0;
    391: T0 = 8'h0;
    default: begin
      T0 = 8'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T5 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T6 = reset ? 1'h0 : restartRegs_0;
  assign T7 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 8'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryStreamer_0(input clk, input reset,
    input  io_restart,
    output[15:0] io_weights_31,
    output[15:0] io_weights_30,
    output[15:0] io_weights_29,
    output[15:0] io_weights_28,
    output[15:0] io_weights_27,
    output[15:0] io_weights_26,
    output[15:0] io_weights_25,
    output[15:0] io_weights_24,
    output[15:0] io_weights_23,
    output[15:0] io_weights_22,
    output[15:0] io_weights_21,
    output[15:0] io_weights_20,
    output[15:0] io_weights_19,
    output[15:0] io_weights_18,
    output[15:0] io_weights_17,
    output[15:0] io_weights_16,
    output[15:0] io_weights_15,
    output[15:0] io_weights_14,
    output[15:0] io_weights_13,
    output[15:0] io_weights_12,
    output[15:0] io_weights_11,
    output[15:0] io_weights_10,
    output[15:0] io_weights_9,
    output[15:0] io_weights_8,
    output[15:0] io_weights_7,
    output[15:0] io_weights_6,
    output[15:0] io_weights_5,
    output[15:0] io_weights_4,
    output[15:0] io_weights_3,
    output[15:0] io_weights_2,
    output[15:0] io_weights_1,
    output[15:0] io_weights_0,
    output[7:0] io_bias
);

  wire[7:0] T34;
  wire[8:0] T0;
  wire[8:0] T1;
  wire[15:0] T2;
  wire[15:0] T3;
  wire[15:0] T4;
  wire[15:0] T5;
  wire[15:0] T6;
  wire[15:0] T7;
  wire[15:0] T8;
  wire[15:0] T9;
  wire[15:0] T10;
  wire[15:0] T11;
  wire[15:0] T12;
  wire[15:0] T13;
  wire[15:0] T14;
  wire[15:0] T15;
  wire[15:0] T16;
  wire[15:0] T17;
  wire[15:0] T18;
  wire[15:0] T19;
  wire[15:0] T20;
  wire[15:0] T21;
  wire[15:0] T22;
  wire[15:0] T23;
  wire[15:0] T24;
  wire[15:0] T25;
  wire[15:0] T26;
  wire[15:0] T27;
  wire[15:0] T28;
  wire[15:0] T29;
  wire[15:0] T30;
  wire[15:0] T31;
  wire[15:0] T32;
  wire[15:0] T33;
  wire MemoryUnit_io_restartOut;
  wire[31:0] MemoryUnit_io_weights;
  wire MemoryUnit_1_io_restartOut;
  wire[31:0] MemoryUnit_1_io_weights;
  wire MemoryUnit_2_io_restartOut;
  wire[31:0] MemoryUnit_2_io_weights;
  wire MemoryUnit_3_io_restartOut;
  wire[31:0] MemoryUnit_3_io_weights;
  wire MemoryUnit_4_io_restartOut;
  wire[31:0] MemoryUnit_4_io_weights;
  wire MemoryUnit_5_io_restartOut;
  wire[31:0] MemoryUnit_5_io_weights;
  wire MemoryUnit_6_io_restartOut;
  wire[31:0] MemoryUnit_6_io_weights;
  wire MemoryUnit_7_io_restartOut;
  wire[31:0] MemoryUnit_7_io_weights;
  wire MemoryUnit_8_io_restartOut;
  wire[31:0] MemoryUnit_8_io_weights;
  wire MemoryUnit_9_io_restartOut;
  wire[31:0] MemoryUnit_9_io_weights;
  wire MemoryUnit_10_io_restartOut;
  wire[31:0] MemoryUnit_10_io_weights;
  wire MemoryUnit_11_io_restartOut;
  wire[31:0] MemoryUnit_11_io_weights;
  wire MemoryUnit_12_io_restartOut;
  wire[31:0] MemoryUnit_12_io_weights;
  wire MemoryUnit_13_io_restartOut;
  wire[31:0] MemoryUnit_13_io_weights;
  wire MemoryUnit_14_io_restartOut;
  wire[31:0] MemoryUnit_14_io_weights;
  wire[31:0] MemoryUnit_15_io_weights;
  wire[7:0] biasMemoryUnit_io_weights;


  assign io_bias = T34;
  assign T34 = T0[7:0];
  assign T0 = T1;
  assign T1 = {1'h0, biasMemoryUnit_io_weights};
  assign io_weights_0 = T2;
  assign T2 = MemoryUnit_io_weights[15:0];
  assign io_weights_1 = T3;
  assign T3 = MemoryUnit_io_weights[31:16];
  assign io_weights_2 = T4;
  assign T4 = MemoryUnit_1_io_weights[15:0];
  assign io_weights_3 = T5;
  assign T5 = MemoryUnit_1_io_weights[31:16];
  assign io_weights_4 = T6;
  assign T6 = MemoryUnit_2_io_weights[15:0];
  assign io_weights_5 = T7;
  assign T7 = MemoryUnit_2_io_weights[31:16];
  assign io_weights_6 = T8;
  assign T8 = MemoryUnit_3_io_weights[15:0];
  assign io_weights_7 = T9;
  assign T9 = MemoryUnit_3_io_weights[31:16];
  assign io_weights_8 = T10;
  assign T10 = MemoryUnit_4_io_weights[15:0];
  assign io_weights_9 = T11;
  assign T11 = MemoryUnit_4_io_weights[31:16];
  assign io_weights_10 = T12;
  assign T12 = MemoryUnit_5_io_weights[15:0];
  assign io_weights_11 = T13;
  assign T13 = MemoryUnit_5_io_weights[31:16];
  assign io_weights_12 = T14;
  assign T14 = MemoryUnit_6_io_weights[15:0];
  assign io_weights_13 = T15;
  assign T15 = MemoryUnit_6_io_weights[31:16];
  assign io_weights_14 = T16;
  assign T16 = MemoryUnit_7_io_weights[15:0];
  assign io_weights_15 = T17;
  assign T17 = MemoryUnit_7_io_weights[31:16];
  assign io_weights_16 = T18;
  assign T18 = MemoryUnit_8_io_weights[15:0];
  assign io_weights_17 = T19;
  assign T19 = MemoryUnit_8_io_weights[31:16];
  assign io_weights_18 = T20;
  assign T20 = MemoryUnit_9_io_weights[15:0];
  assign io_weights_19 = T21;
  assign T21 = MemoryUnit_9_io_weights[31:16];
  assign io_weights_20 = T22;
  assign T22 = MemoryUnit_10_io_weights[15:0];
  assign io_weights_21 = T23;
  assign T23 = MemoryUnit_10_io_weights[31:16];
  assign io_weights_22 = T24;
  assign T24 = MemoryUnit_11_io_weights[15:0];
  assign io_weights_23 = T25;
  assign T25 = MemoryUnit_11_io_weights[31:16];
  assign io_weights_24 = T26;
  assign T26 = MemoryUnit_12_io_weights[15:0];
  assign io_weights_25 = T27;
  assign T27 = MemoryUnit_12_io_weights[31:16];
  assign io_weights_26 = T28;
  assign T28 = MemoryUnit_13_io_weights[15:0];
  assign io_weights_27 = T29;
  assign T29 = MemoryUnit_13_io_weights[31:16];
  assign io_weights_28 = T30;
  assign T30 = MemoryUnit_14_io_weights[15:0];
  assign io_weights_29 = T31;
  assign T31 = MemoryUnit_14_io_weights[31:16];
  assign io_weights_30 = T32;
  assign T32 = MemoryUnit_15_io_weights[15:0];
  assign io_weights_31 = T33;
  assign T33 = MemoryUnit_15_io_weights[31:16];
  MemoryUnit_0 MemoryUnit(.clk(clk), .reset(reset),
       .io_restartIn( io_restart ),
       .io_restartOut( MemoryUnit_io_restartOut ),
       .io_weights( MemoryUnit_io_weights )
  );
  MemoryUnit_1 MemoryUnit_1(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_io_restartOut ),
       .io_restartOut( MemoryUnit_1_io_restartOut ),
       .io_weights( MemoryUnit_1_io_weights )
  );
  MemoryUnit_2 MemoryUnit_2(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_1_io_restartOut ),
       .io_restartOut( MemoryUnit_2_io_restartOut ),
       .io_weights( MemoryUnit_2_io_weights )
  );
  MemoryUnit_3 MemoryUnit_3(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_2_io_restartOut ),
       .io_restartOut( MemoryUnit_3_io_restartOut ),
       .io_weights( MemoryUnit_3_io_weights )
  );
  MemoryUnit_4 MemoryUnit_4(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_3_io_restartOut ),
       .io_restartOut( MemoryUnit_4_io_restartOut ),
       .io_weights( MemoryUnit_4_io_weights )
  );
  MemoryUnit_5 MemoryUnit_5(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_4_io_restartOut ),
       .io_restartOut( MemoryUnit_5_io_restartOut ),
       .io_weights( MemoryUnit_5_io_weights )
  );
  MemoryUnit_6 MemoryUnit_6(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_5_io_restartOut ),
       .io_restartOut( MemoryUnit_6_io_restartOut ),
       .io_weights( MemoryUnit_6_io_weights )
  );
  MemoryUnit_7 MemoryUnit_7(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_6_io_restartOut ),
       .io_restartOut( MemoryUnit_7_io_restartOut ),
       .io_weights( MemoryUnit_7_io_weights )
  );
  MemoryUnit_8 MemoryUnit_8(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_7_io_restartOut ),
       .io_restartOut( MemoryUnit_8_io_restartOut ),
       .io_weights( MemoryUnit_8_io_weights )
  );
  MemoryUnit_9 MemoryUnit_9(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_8_io_restartOut ),
       .io_restartOut( MemoryUnit_9_io_restartOut ),
       .io_weights( MemoryUnit_9_io_weights )
  );
  MemoryUnit_10 MemoryUnit_10(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_9_io_restartOut ),
       .io_restartOut( MemoryUnit_10_io_restartOut ),
       .io_weights( MemoryUnit_10_io_weights )
  );
  MemoryUnit_11 MemoryUnit_11(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_10_io_restartOut ),
       .io_restartOut( MemoryUnit_11_io_restartOut ),
       .io_weights( MemoryUnit_11_io_weights )
  );
  MemoryUnit_12 MemoryUnit_12(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_11_io_restartOut ),
       .io_restartOut( MemoryUnit_12_io_restartOut ),
       .io_weights( MemoryUnit_12_io_weights )
  );
  MemoryUnit_13 MemoryUnit_13(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_12_io_restartOut ),
       .io_restartOut( MemoryUnit_13_io_restartOut ),
       .io_weights( MemoryUnit_13_io_weights )
  );
  MemoryUnit_14 MemoryUnit_14(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_13_io_restartOut ),
       .io_restartOut( MemoryUnit_14_io_restartOut ),
       .io_weights( MemoryUnit_14_io_weights )
  );
  MemoryUnit_15 MemoryUnit_15(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_14_io_restartOut ),
       //.io_restartOut(  )
       .io_weights( MemoryUnit_15_io_weights )
  );
  MemoryUnit_16 biasMemoryUnit(.clk(clk), .reset(reset),
       .io_restartIn( io_restart ),
       //.io_restartOut(  )
       .io_weights( biasMemoryUnit_io_weights )
  );
endmodule

module Warp_0(input clk, input reset,
    input [15:0] io_xIn_3,
    input [15:0] io_xIn_2,
    input [15:0] io_xIn_1,
    input [15:0] io_xIn_0,
    input  io_start,
    output io_ready,
    output io_startOut,
    output io_xOut_3,
    output io_xOut_2,
    output io_xOut_1,
    output io_xOut_0,
    output io_xOutValid,
    input  io_pipeReady,
    output io_done
);

  wire[9:0] T508;
  wire[10:0] T0;
  wire[10:0] T1;
  wire[9:0] T509;
  wire[10:0] T2;
  wire[10:0] T3;
  wire[9:0] T510;
  wire[10:0] T4;
  wire[10:0] T5;
  wire[9:0] T511;
  wire[10:0] T6;
  wire[10:0] T7;
  wire[9:0] T512;
  wire[10:0] T8;
  wire[10:0] T9;
  wire[9:0] T513;
  wire[10:0] T10;
  wire[10:0] T11;
  wire[9:0] T514;
  wire[10:0] T12;
  wire[10:0] T13;
  wire[9:0] T515;
  wire[10:0] T14;
  wire[10:0] T15;
  wire[9:0] T516;
  wire[10:0] T16;
  wire[10:0] T17;
  wire[9:0] T517;
  wire[10:0] T18;
  wire[10:0] T19;
  wire[9:0] T518;
  wire[10:0] T20;
  wire[10:0] T21;
  wire[9:0] T519;
  wire[10:0] T22;
  wire[10:0] T23;
  wire[9:0] T520;
  wire[10:0] T24;
  wire[10:0] T25;
  wire[9:0] T521;
  wire[10:0] T26;
  wire[10:0] T27;
  wire[9:0] T522;
  wire[10:0] T28;
  wire[10:0] T29;
  wire[9:0] T523;
  wire[10:0] T30;
  wire[10:0] T31;
  wire[9:0] T524;
  wire[10:0] T32;
  wire[10:0] T33;
  wire[9:0] T525;
  wire[10:0] T34;
  wire[10:0] T35;
  wire[9:0] T526;
  wire[10:0] T36;
  wire[10:0] T37;
  wire[9:0] T527;
  wire[10:0] T38;
  wire[10:0] T39;
  wire[9:0] T528;
  wire[10:0] T40;
  wire[10:0] T41;
  wire[9:0] T529;
  wire[10:0] T42;
  wire[10:0] T43;
  wire[9:0] T530;
  wire[10:0] T44;
  wire[10:0] T45;
  wire[9:0] T531;
  wire[10:0] T46;
  wire[10:0] T47;
  wire[9:0] T532;
  wire[10:0] T48;
  wire[10:0] T49;
  wire[9:0] T533;
  wire[10:0] T50;
  wire[10:0] T51;
  wire[9:0] T534;
  wire[10:0] T52;
  wire[10:0] T53;
  wire[9:0] T535;
  wire[10:0] T54;
  wire[10:0] T55;
  wire[9:0] T536;
  wire[10:0] T56;
  wire[10:0] T57;
  wire[9:0] T537;
  wire[10:0] T58;
  wire[10:0] T59;
  wire[9:0] T538;
  wire[10:0] T60;
  wire[10:0] T61;
  wire[9:0] T539;
  wire[10:0] T62;
  wire[10:0] T63;
  wire[9:0] T540;
  wire[10:0] T64;
  wire[10:0] T65;
  wire[9:0] T541;
  wire[10:0] T66;
  wire[10:0] T67;
  wire[9:0] T542;
  wire[10:0] T68;
  wire[10:0] T69;
  wire[9:0] T543;
  wire[10:0] T70;
  wire[10:0] T71;
  wire[9:0] T544;
  wire[10:0] T72;
  wire[10:0] T73;
  wire[9:0] T545;
  wire[10:0] T74;
  wire[10:0] T75;
  wire[9:0] T546;
  wire[10:0] T76;
  wire[10:0] T77;
  wire[9:0] T547;
  wire[10:0] T78;
  wire[10:0] T79;
  wire[9:0] T548;
  wire[10:0] T80;
  wire[10:0] T81;
  wire[9:0] T549;
  wire[10:0] T82;
  wire[10:0] T83;
  wire[9:0] T550;
  wire[10:0] T84;
  wire[10:0] T85;
  wire[9:0] T551;
  wire[10:0] T86;
  wire[10:0] T87;
  wire[9:0] T552;
  wire[10:0] T88;
  wire[10:0] T89;
  wire[9:0] T553;
  wire[10:0] T90;
  wire[10:0] T91;
  wire[9:0] T554;
  wire[10:0] T92;
  wire[10:0] T93;
  wire[9:0] T555;
  wire[10:0] T94;
  wire[10:0] T95;
  wire[9:0] T556;
  wire[10:0] T96;
  wire[10:0] T97;
  wire[9:0] T557;
  wire[10:0] T98;
  wire[10:0] T99;
  wire[9:0] T558;
  wire[10:0] T100;
  wire[10:0] T101;
  wire[9:0] T559;
  wire[10:0] T102;
  wire[10:0] T103;
  wire[9:0] T560;
  wire[10:0] T104;
  wire[10:0] T105;
  wire[9:0] T561;
  wire[10:0] T106;
  wire[10:0] T107;
  wire[9:0] T562;
  wire[10:0] T108;
  wire[10:0] T109;
  wire[9:0] T563;
  wire[10:0] T110;
  wire[10:0] T111;
  wire[9:0] T564;
  wire[10:0] T112;
  wire[10:0] T113;
  wire[9:0] T565;
  wire[10:0] T114;
  wire[10:0] T115;
  wire[9:0] T566;
  wire[10:0] T116;
  wire[10:0] T117;
  wire[9:0] T567;
  wire[10:0] T118;
  wire[10:0] T119;
  wire[9:0] T568;
  wire[10:0] T120;
  wire[10:0] T121;
  wire[9:0] T569;
  wire[10:0] T122;
  wire[10:0] T123;
  wire[9:0] T570;
  wire[10:0] T124;
  wire[10:0] T125;
  wire[9:0] T571;
  wire[10:0] T126;
  wire[10:0] T127;
  wire[9:0] T572;
  wire[10:0] T128;
  wire[10:0] T129;
  wire[9:0] T573;
  wire[10:0] T130;
  wire[10:0] T131;
  wire[9:0] T574;
  wire[10:0] T132;
  wire[10:0] T133;
  wire[9:0] T575;
  wire[10:0] T134;
  wire[10:0] T135;
  wire[9:0] T576;
  wire[10:0] T136;
  wire[10:0] T137;
  wire[9:0] T577;
  wire[10:0] T138;
  wire[10:0] T139;
  wire[9:0] T578;
  wire[10:0] T140;
  wire[10:0] T141;
  wire[9:0] T579;
  wire[10:0] T142;
  wire[10:0] T143;
  wire[9:0] T580;
  wire[10:0] T144;
  wire[10:0] T145;
  wire[9:0] T581;
  wire[10:0] T146;
  wire[10:0] T147;
  wire[9:0] T582;
  wire[10:0] T148;
  wire[10:0] T149;
  wire[9:0] T583;
  wire[10:0] T150;
  wire[10:0] T151;
  wire[9:0] T584;
  wire[10:0] T152;
  wire[10:0] T153;
  wire[9:0] T585;
  wire[10:0] T154;
  wire[10:0] T155;
  wire[9:0] T586;
  wire[10:0] T156;
  wire[10:0] T157;
  wire[9:0] T587;
  wire[10:0] T158;
  wire[10:0] T159;
  wire[9:0] T588;
  wire[10:0] T160;
  wire[10:0] T161;
  wire[9:0] T589;
  wire[10:0] T162;
  wire[10:0] T163;
  wire[9:0] T590;
  wire[10:0] T164;
  wire[10:0] T165;
  wire[9:0] T591;
  wire[10:0] T166;
  wire[10:0] T167;
  wire[9:0] T592;
  wire[10:0] T168;
  wire[10:0] T169;
  wire[9:0] T593;
  wire[10:0] T170;
  wire[10:0] T171;
  wire[9:0] T594;
  wire[10:0] T172;
  wire[10:0] T173;
  wire[9:0] T595;
  wire[10:0] T174;
  wire[10:0] T175;
  wire[9:0] T596;
  wire[10:0] T176;
  wire[10:0] T177;
  wire[9:0] T597;
  wire[10:0] T178;
  wire[10:0] T179;
  wire[9:0] T598;
  wire[10:0] T180;
  wire[10:0] T181;
  wire[9:0] T599;
  wire[10:0] T182;
  wire[10:0] T183;
  wire[9:0] T600;
  wire[10:0] T184;
  wire[10:0] T185;
  wire[9:0] T601;
  wire[10:0] T186;
  wire[10:0] T187;
  wire[9:0] T602;
  wire[10:0] T188;
  wire[10:0] T189;
  wire[9:0] T603;
  wire[10:0] T190;
  wire[10:0] T191;
  wire[9:0] T604;
  wire[10:0] T192;
  wire[10:0] T193;
  wire[9:0] T605;
  wire[10:0] T194;
  wire[10:0] T195;
  wire[9:0] T606;
  wire[10:0] T196;
  wire[10:0] T197;
  wire[9:0] T607;
  wire[10:0] T198;
  wire[10:0] T199;
  wire[9:0] T608;
  wire[10:0] T200;
  wire[10:0] T201;
  wire[9:0] T609;
  wire[10:0] T202;
  wire[10:0] T203;
  wire[9:0] T610;
  wire[10:0] T204;
  wire[10:0] T205;
  wire[9:0] T611;
  wire[10:0] T206;
  wire[10:0] T207;
  wire[9:0] T612;
  wire[10:0] T208;
  wire[10:0] T209;
  wire[9:0] T613;
  wire[10:0] T210;
  wire[10:0] T211;
  wire[9:0] T614;
  wire[10:0] T212;
  wire[10:0] T213;
  wire[9:0] T615;
  wire[10:0] T214;
  wire[10:0] T215;
  wire[9:0] T616;
  wire[10:0] T216;
  wire[10:0] T217;
  wire[9:0] T617;
  wire[10:0] T218;
  wire[10:0] T219;
  wire[9:0] T618;
  wire[10:0] T220;
  wire[10:0] T221;
  wire[9:0] T619;
  wire[10:0] T222;
  wire[10:0] T223;
  wire[9:0] T620;
  wire[10:0] T224;
  wire[10:0] T225;
  wire[9:0] T621;
  wire[10:0] T226;
  wire[10:0] T227;
  wire[9:0] T622;
  wire[10:0] T228;
  wire[10:0] T229;
  wire[9:0] T623;
  wire[10:0] T230;
  wire[10:0] T231;
  wire[9:0] T624;
  wire[10:0] T232;
  wire[10:0] T233;
  wire[9:0] T625;
  wire[10:0] T234;
  wire[10:0] T235;
  wire[9:0] T626;
  wire[10:0] T236;
  wire[10:0] T237;
  wire[9:0] T627;
  wire[10:0] T238;
  wire[10:0] T239;
  wire[9:0] T628;
  wire[10:0] T240;
  wire[10:0] T241;
  wire[9:0] T629;
  wire[10:0] T242;
  wire[10:0] T243;
  wire[9:0] T630;
  wire[10:0] T244;
  wire[10:0] T245;
  wire[9:0] T631;
  wire[10:0] T246;
  wire[10:0] T247;
  wire[9:0] T632;
  wire[10:0] T248;
  wire[10:0] T249;
  wire[9:0] T633;
  wire[10:0] T250;
  wire[10:0] T251;
  wire[9:0] T634;
  wire[10:0] T252;
  wire[10:0] T253;
  wire[9:0] T635;
  wire[10:0] T254;
  wire[10:0] T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire[4:0] T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire[4:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire[4:0] T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire[4:0] T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire T492;
  wire T493;
  wire T494;
  wire T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;
  wire T500;
  wire T501;
  wire T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire Activation_io_out_31;
  wire Activation_io_out_30;
  wire Activation_io_out_29;
  wire Activation_io_out_28;
  wire Activation_io_out_27;
  wire Activation_io_out_26;
  wire Activation_io_out_25;
  wire Activation_io_out_24;
  wire Activation_io_out_23;
  wire Activation_io_out_22;
  wire Activation_io_out_21;
  wire Activation_io_out_20;
  wire Activation_io_out_19;
  wire Activation_io_out_18;
  wire Activation_io_out_17;
  wire Activation_io_out_16;
  wire Activation_io_out_15;
  wire Activation_io_out_14;
  wire Activation_io_out_13;
  wire Activation_io_out_12;
  wire Activation_io_out_11;
  wire Activation_io_out_10;
  wire Activation_io_out_9;
  wire Activation_io_out_8;
  wire Activation_io_out_7;
  wire Activation_io_out_6;
  wire Activation_io_out_5;
  wire Activation_io_out_4;
  wire Activation_io_out_3;
  wire Activation_io_out_2;
  wire Activation_io_out_1;
  wire Activation_io_out_0;
  wire Activation_1_io_out_31;
  wire Activation_1_io_out_30;
  wire Activation_1_io_out_29;
  wire Activation_1_io_out_28;
  wire Activation_1_io_out_27;
  wire Activation_1_io_out_26;
  wire Activation_1_io_out_25;
  wire Activation_1_io_out_24;
  wire Activation_1_io_out_23;
  wire Activation_1_io_out_22;
  wire Activation_1_io_out_21;
  wire Activation_1_io_out_20;
  wire Activation_1_io_out_19;
  wire Activation_1_io_out_18;
  wire Activation_1_io_out_17;
  wire Activation_1_io_out_16;
  wire Activation_1_io_out_15;
  wire Activation_1_io_out_14;
  wire Activation_1_io_out_13;
  wire Activation_1_io_out_12;
  wire Activation_1_io_out_11;
  wire Activation_1_io_out_10;
  wire Activation_1_io_out_9;
  wire Activation_1_io_out_8;
  wire Activation_1_io_out_7;
  wire Activation_1_io_out_6;
  wire Activation_1_io_out_5;
  wire Activation_1_io_out_4;
  wire Activation_1_io_out_3;
  wire Activation_1_io_out_2;
  wire Activation_1_io_out_1;
  wire Activation_1_io_out_0;
  wire Activation_2_io_out_31;
  wire Activation_2_io_out_30;
  wire Activation_2_io_out_29;
  wire Activation_2_io_out_28;
  wire Activation_2_io_out_27;
  wire Activation_2_io_out_26;
  wire Activation_2_io_out_25;
  wire Activation_2_io_out_24;
  wire Activation_2_io_out_23;
  wire Activation_2_io_out_22;
  wire Activation_2_io_out_21;
  wire Activation_2_io_out_20;
  wire Activation_2_io_out_19;
  wire Activation_2_io_out_18;
  wire Activation_2_io_out_17;
  wire Activation_2_io_out_16;
  wire Activation_2_io_out_15;
  wire Activation_2_io_out_14;
  wire Activation_2_io_out_13;
  wire Activation_2_io_out_12;
  wire Activation_2_io_out_11;
  wire Activation_2_io_out_10;
  wire Activation_2_io_out_9;
  wire Activation_2_io_out_8;
  wire Activation_2_io_out_7;
  wire Activation_2_io_out_6;
  wire Activation_2_io_out_5;
  wire Activation_2_io_out_4;
  wire Activation_2_io_out_3;
  wire Activation_2_io_out_2;
  wire Activation_2_io_out_1;
  wire Activation_2_io_out_0;
  wire Activation_3_io_out_31;
  wire Activation_3_io_out_30;
  wire Activation_3_io_out_29;
  wire Activation_3_io_out_28;
  wire Activation_3_io_out_27;
  wire Activation_3_io_out_26;
  wire Activation_3_io_out_25;
  wire Activation_3_io_out_24;
  wire Activation_3_io_out_23;
  wire Activation_3_io_out_22;
  wire Activation_3_io_out_21;
  wire Activation_3_io_out_20;
  wire Activation_3_io_out_19;
  wire Activation_3_io_out_18;
  wire Activation_3_io_out_17;
  wire Activation_3_io_out_16;
  wire Activation_3_io_out_15;
  wire Activation_3_io_out_14;
  wire Activation_3_io_out_13;
  wire Activation_3_io_out_12;
  wire Activation_3_io_out_11;
  wire Activation_3_io_out_10;
  wire Activation_3_io_out_9;
  wire Activation_3_io_out_8;
  wire Activation_3_io_out_7;
  wire Activation_3_io_out_6;
  wire Activation_3_io_out_5;
  wire Activation_3_io_out_4;
  wire Activation_3_io_out_3;
  wire Activation_3_io_out_2;
  wire Activation_3_io_out_1;
  wire Activation_3_io_out_0;
  wire control_io_ready;
  wire control_io_valid;
  wire control_io_done;
  wire[4:0] control_io_selectX;
  wire control_io_memoryRestart;
  wire control_io_chainRestart;
  wire[9:0] Chain_io_ys_31;
  wire[9:0] Chain_io_ys_30;
  wire[9:0] Chain_io_ys_29;
  wire[9:0] Chain_io_ys_28;
  wire[9:0] Chain_io_ys_27;
  wire[9:0] Chain_io_ys_26;
  wire[9:0] Chain_io_ys_25;
  wire[9:0] Chain_io_ys_24;
  wire[9:0] Chain_io_ys_23;
  wire[9:0] Chain_io_ys_22;
  wire[9:0] Chain_io_ys_21;
  wire[9:0] Chain_io_ys_20;
  wire[9:0] Chain_io_ys_19;
  wire[9:0] Chain_io_ys_18;
  wire[9:0] Chain_io_ys_17;
  wire[9:0] Chain_io_ys_16;
  wire[9:0] Chain_io_ys_15;
  wire[9:0] Chain_io_ys_14;
  wire[9:0] Chain_io_ys_13;
  wire[9:0] Chain_io_ys_12;
  wire[9:0] Chain_io_ys_11;
  wire[9:0] Chain_io_ys_10;
  wire[9:0] Chain_io_ys_9;
  wire[9:0] Chain_io_ys_8;
  wire[9:0] Chain_io_ys_7;
  wire[9:0] Chain_io_ys_6;
  wire[9:0] Chain_io_ys_5;
  wire[9:0] Chain_io_ys_4;
  wire[9:0] Chain_io_ys_3;
  wire[9:0] Chain_io_ys_2;
  wire[9:0] Chain_io_ys_1;
  wire[9:0] Chain_io_ys_0;
  wire[9:0] Chain_1_io_ys_31;
  wire[9:0] Chain_1_io_ys_30;
  wire[9:0] Chain_1_io_ys_29;
  wire[9:0] Chain_1_io_ys_28;
  wire[9:0] Chain_1_io_ys_27;
  wire[9:0] Chain_1_io_ys_26;
  wire[9:0] Chain_1_io_ys_25;
  wire[9:0] Chain_1_io_ys_24;
  wire[9:0] Chain_1_io_ys_23;
  wire[9:0] Chain_1_io_ys_22;
  wire[9:0] Chain_1_io_ys_21;
  wire[9:0] Chain_1_io_ys_20;
  wire[9:0] Chain_1_io_ys_19;
  wire[9:0] Chain_1_io_ys_18;
  wire[9:0] Chain_1_io_ys_17;
  wire[9:0] Chain_1_io_ys_16;
  wire[9:0] Chain_1_io_ys_15;
  wire[9:0] Chain_1_io_ys_14;
  wire[9:0] Chain_1_io_ys_13;
  wire[9:0] Chain_1_io_ys_12;
  wire[9:0] Chain_1_io_ys_11;
  wire[9:0] Chain_1_io_ys_10;
  wire[9:0] Chain_1_io_ys_9;
  wire[9:0] Chain_1_io_ys_8;
  wire[9:0] Chain_1_io_ys_7;
  wire[9:0] Chain_1_io_ys_6;
  wire[9:0] Chain_1_io_ys_5;
  wire[9:0] Chain_1_io_ys_4;
  wire[9:0] Chain_1_io_ys_3;
  wire[9:0] Chain_1_io_ys_2;
  wire[9:0] Chain_1_io_ys_1;
  wire[9:0] Chain_1_io_ys_0;
  wire[9:0] Chain_2_io_ys_31;
  wire[9:0] Chain_2_io_ys_30;
  wire[9:0] Chain_2_io_ys_29;
  wire[9:0] Chain_2_io_ys_28;
  wire[9:0] Chain_2_io_ys_27;
  wire[9:0] Chain_2_io_ys_26;
  wire[9:0] Chain_2_io_ys_25;
  wire[9:0] Chain_2_io_ys_24;
  wire[9:0] Chain_2_io_ys_23;
  wire[9:0] Chain_2_io_ys_22;
  wire[9:0] Chain_2_io_ys_21;
  wire[9:0] Chain_2_io_ys_20;
  wire[9:0] Chain_2_io_ys_19;
  wire[9:0] Chain_2_io_ys_18;
  wire[9:0] Chain_2_io_ys_17;
  wire[9:0] Chain_2_io_ys_16;
  wire[9:0] Chain_2_io_ys_15;
  wire[9:0] Chain_2_io_ys_14;
  wire[9:0] Chain_2_io_ys_13;
  wire[9:0] Chain_2_io_ys_12;
  wire[9:0] Chain_2_io_ys_11;
  wire[9:0] Chain_2_io_ys_10;
  wire[9:0] Chain_2_io_ys_9;
  wire[9:0] Chain_2_io_ys_8;
  wire[9:0] Chain_2_io_ys_7;
  wire[9:0] Chain_2_io_ys_6;
  wire[9:0] Chain_2_io_ys_5;
  wire[9:0] Chain_2_io_ys_4;
  wire[9:0] Chain_2_io_ys_3;
  wire[9:0] Chain_2_io_ys_2;
  wire[9:0] Chain_2_io_ys_1;
  wire[9:0] Chain_2_io_ys_0;
  wire[9:0] Chain_3_io_ys_31;
  wire[9:0] Chain_3_io_ys_30;
  wire[9:0] Chain_3_io_ys_29;
  wire[9:0] Chain_3_io_ys_28;
  wire[9:0] Chain_3_io_ys_27;
  wire[9:0] Chain_3_io_ys_26;
  wire[9:0] Chain_3_io_ys_25;
  wire[9:0] Chain_3_io_ys_24;
  wire[9:0] Chain_3_io_ys_23;
  wire[9:0] Chain_3_io_ys_22;
  wire[9:0] Chain_3_io_ys_21;
  wire[9:0] Chain_3_io_ys_20;
  wire[9:0] Chain_3_io_ys_19;
  wire[9:0] Chain_3_io_ys_18;
  wire[9:0] Chain_3_io_ys_17;
  wire[9:0] Chain_3_io_ys_16;
  wire[9:0] Chain_3_io_ys_15;
  wire[9:0] Chain_3_io_ys_14;
  wire[9:0] Chain_3_io_ys_13;
  wire[9:0] Chain_3_io_ys_12;
  wire[9:0] Chain_3_io_ys_11;
  wire[9:0] Chain_3_io_ys_10;
  wire[9:0] Chain_3_io_ys_9;
  wire[9:0] Chain_3_io_ys_8;
  wire[9:0] Chain_3_io_ys_7;
  wire[9:0] Chain_3_io_ys_6;
  wire[9:0] Chain_3_io_ys_5;
  wire[9:0] Chain_3_io_ys_4;
  wire[9:0] Chain_3_io_ys_3;
  wire[9:0] Chain_3_io_ys_2;
  wire[9:0] Chain_3_io_ys_1;
  wire[9:0] Chain_3_io_ys_0;
  wire[15:0] memoryStreamer_io_weights_31;
  wire[15:0] memoryStreamer_io_weights_30;
  wire[15:0] memoryStreamer_io_weights_29;
  wire[15:0] memoryStreamer_io_weights_28;
  wire[15:0] memoryStreamer_io_weights_27;
  wire[15:0] memoryStreamer_io_weights_26;
  wire[15:0] memoryStreamer_io_weights_25;
  wire[15:0] memoryStreamer_io_weights_24;
  wire[15:0] memoryStreamer_io_weights_23;
  wire[15:0] memoryStreamer_io_weights_22;
  wire[15:0] memoryStreamer_io_weights_21;
  wire[15:0] memoryStreamer_io_weights_20;
  wire[15:0] memoryStreamer_io_weights_19;
  wire[15:0] memoryStreamer_io_weights_18;
  wire[15:0] memoryStreamer_io_weights_17;
  wire[15:0] memoryStreamer_io_weights_16;
  wire[15:0] memoryStreamer_io_weights_15;
  wire[15:0] memoryStreamer_io_weights_14;
  wire[15:0] memoryStreamer_io_weights_13;
  wire[15:0] memoryStreamer_io_weights_12;
  wire[15:0] memoryStreamer_io_weights_11;
  wire[15:0] memoryStreamer_io_weights_10;
  wire[15:0] memoryStreamer_io_weights_9;
  wire[15:0] memoryStreamer_io_weights_8;
  wire[15:0] memoryStreamer_io_weights_7;
  wire[15:0] memoryStreamer_io_weights_6;
  wire[15:0] memoryStreamer_io_weights_5;
  wire[15:0] memoryStreamer_io_weights_4;
  wire[15:0] memoryStreamer_io_weights_3;
  wire[15:0] memoryStreamer_io_weights_2;
  wire[15:0] memoryStreamer_io_weights_1;
  wire[15:0] memoryStreamer_io_weights_0;
  wire[7:0] memoryStreamer_io_bias;


  assign T508 = T0[9:0];
  assign T0 = T1;
  assign T1 = {1'h0, Chain_3_io_ys_0};
  assign T509 = T2[9:0];
  assign T2 = T3;
  assign T3 = {1'h0, Chain_3_io_ys_1};
  assign T510 = T4[9:0];
  assign T4 = T5;
  assign T5 = {1'h0, Chain_3_io_ys_2};
  assign T511 = T6[9:0];
  assign T6 = T7;
  assign T7 = {1'h0, Chain_3_io_ys_3};
  assign T512 = T8[9:0];
  assign T8 = T9;
  assign T9 = {1'h0, Chain_3_io_ys_4};
  assign T513 = T10[9:0];
  assign T10 = T11;
  assign T11 = {1'h0, Chain_3_io_ys_5};
  assign T514 = T12[9:0];
  assign T12 = T13;
  assign T13 = {1'h0, Chain_3_io_ys_6};
  assign T515 = T14[9:0];
  assign T14 = T15;
  assign T15 = {1'h0, Chain_3_io_ys_7};
  assign T516 = T16[9:0];
  assign T16 = T17;
  assign T17 = {1'h0, Chain_3_io_ys_8};
  assign T517 = T18[9:0];
  assign T18 = T19;
  assign T19 = {1'h0, Chain_3_io_ys_9};
  assign T518 = T20[9:0];
  assign T20 = T21;
  assign T21 = {1'h0, Chain_3_io_ys_10};
  assign T519 = T22[9:0];
  assign T22 = T23;
  assign T23 = {1'h0, Chain_3_io_ys_11};
  assign T520 = T24[9:0];
  assign T24 = T25;
  assign T25 = {1'h0, Chain_3_io_ys_12};
  assign T521 = T26[9:0];
  assign T26 = T27;
  assign T27 = {1'h0, Chain_3_io_ys_13};
  assign T522 = T28[9:0];
  assign T28 = T29;
  assign T29 = {1'h0, Chain_3_io_ys_14};
  assign T523 = T30[9:0];
  assign T30 = T31;
  assign T31 = {1'h0, Chain_3_io_ys_15};
  assign T524 = T32[9:0];
  assign T32 = T33;
  assign T33 = {1'h0, Chain_3_io_ys_16};
  assign T525 = T34[9:0];
  assign T34 = T35;
  assign T35 = {1'h0, Chain_3_io_ys_17};
  assign T526 = T36[9:0];
  assign T36 = T37;
  assign T37 = {1'h0, Chain_3_io_ys_18};
  assign T527 = T38[9:0];
  assign T38 = T39;
  assign T39 = {1'h0, Chain_3_io_ys_19};
  assign T528 = T40[9:0];
  assign T40 = T41;
  assign T41 = {1'h0, Chain_3_io_ys_20};
  assign T529 = T42[9:0];
  assign T42 = T43;
  assign T43 = {1'h0, Chain_3_io_ys_21};
  assign T530 = T44[9:0];
  assign T44 = T45;
  assign T45 = {1'h0, Chain_3_io_ys_22};
  assign T531 = T46[9:0];
  assign T46 = T47;
  assign T47 = {1'h0, Chain_3_io_ys_23};
  assign T532 = T48[9:0];
  assign T48 = T49;
  assign T49 = {1'h0, Chain_3_io_ys_24};
  assign T533 = T50[9:0];
  assign T50 = T51;
  assign T51 = {1'h0, Chain_3_io_ys_25};
  assign T534 = T52[9:0];
  assign T52 = T53;
  assign T53 = {1'h0, Chain_3_io_ys_26};
  assign T535 = T54[9:0];
  assign T54 = T55;
  assign T55 = {1'h0, Chain_3_io_ys_27};
  assign T536 = T56[9:0];
  assign T56 = T57;
  assign T57 = {1'h0, Chain_3_io_ys_28};
  assign T537 = T58[9:0];
  assign T58 = T59;
  assign T59 = {1'h0, Chain_3_io_ys_29};
  assign T538 = T60[9:0];
  assign T60 = T61;
  assign T61 = {1'h0, Chain_3_io_ys_30};
  assign T539 = T62[9:0];
  assign T62 = T63;
  assign T63 = {1'h0, Chain_3_io_ys_31};
  assign T540 = T64[9:0];
  assign T64 = T65;
  assign T65 = {1'h0, Chain_2_io_ys_0};
  assign T541 = T66[9:0];
  assign T66 = T67;
  assign T67 = {1'h0, Chain_2_io_ys_1};
  assign T542 = T68[9:0];
  assign T68 = T69;
  assign T69 = {1'h0, Chain_2_io_ys_2};
  assign T543 = T70[9:0];
  assign T70 = T71;
  assign T71 = {1'h0, Chain_2_io_ys_3};
  assign T544 = T72[9:0];
  assign T72 = T73;
  assign T73 = {1'h0, Chain_2_io_ys_4};
  assign T545 = T74[9:0];
  assign T74 = T75;
  assign T75 = {1'h0, Chain_2_io_ys_5};
  assign T546 = T76[9:0];
  assign T76 = T77;
  assign T77 = {1'h0, Chain_2_io_ys_6};
  assign T547 = T78[9:0];
  assign T78 = T79;
  assign T79 = {1'h0, Chain_2_io_ys_7};
  assign T548 = T80[9:0];
  assign T80 = T81;
  assign T81 = {1'h0, Chain_2_io_ys_8};
  assign T549 = T82[9:0];
  assign T82 = T83;
  assign T83 = {1'h0, Chain_2_io_ys_9};
  assign T550 = T84[9:0];
  assign T84 = T85;
  assign T85 = {1'h0, Chain_2_io_ys_10};
  assign T551 = T86[9:0];
  assign T86 = T87;
  assign T87 = {1'h0, Chain_2_io_ys_11};
  assign T552 = T88[9:0];
  assign T88 = T89;
  assign T89 = {1'h0, Chain_2_io_ys_12};
  assign T553 = T90[9:0];
  assign T90 = T91;
  assign T91 = {1'h0, Chain_2_io_ys_13};
  assign T554 = T92[9:0];
  assign T92 = T93;
  assign T93 = {1'h0, Chain_2_io_ys_14};
  assign T555 = T94[9:0];
  assign T94 = T95;
  assign T95 = {1'h0, Chain_2_io_ys_15};
  assign T556 = T96[9:0];
  assign T96 = T97;
  assign T97 = {1'h0, Chain_2_io_ys_16};
  assign T557 = T98[9:0];
  assign T98 = T99;
  assign T99 = {1'h0, Chain_2_io_ys_17};
  assign T558 = T100[9:0];
  assign T100 = T101;
  assign T101 = {1'h0, Chain_2_io_ys_18};
  assign T559 = T102[9:0];
  assign T102 = T103;
  assign T103 = {1'h0, Chain_2_io_ys_19};
  assign T560 = T104[9:0];
  assign T104 = T105;
  assign T105 = {1'h0, Chain_2_io_ys_20};
  assign T561 = T106[9:0];
  assign T106 = T107;
  assign T107 = {1'h0, Chain_2_io_ys_21};
  assign T562 = T108[9:0];
  assign T108 = T109;
  assign T109 = {1'h0, Chain_2_io_ys_22};
  assign T563 = T110[9:0];
  assign T110 = T111;
  assign T111 = {1'h0, Chain_2_io_ys_23};
  assign T564 = T112[9:0];
  assign T112 = T113;
  assign T113 = {1'h0, Chain_2_io_ys_24};
  assign T565 = T114[9:0];
  assign T114 = T115;
  assign T115 = {1'h0, Chain_2_io_ys_25};
  assign T566 = T116[9:0];
  assign T116 = T117;
  assign T117 = {1'h0, Chain_2_io_ys_26};
  assign T567 = T118[9:0];
  assign T118 = T119;
  assign T119 = {1'h0, Chain_2_io_ys_27};
  assign T568 = T120[9:0];
  assign T120 = T121;
  assign T121 = {1'h0, Chain_2_io_ys_28};
  assign T569 = T122[9:0];
  assign T122 = T123;
  assign T123 = {1'h0, Chain_2_io_ys_29};
  assign T570 = T124[9:0];
  assign T124 = T125;
  assign T125 = {1'h0, Chain_2_io_ys_30};
  assign T571 = T126[9:0];
  assign T126 = T127;
  assign T127 = {1'h0, Chain_2_io_ys_31};
  assign T572 = T128[9:0];
  assign T128 = T129;
  assign T129 = {1'h0, Chain_1_io_ys_0};
  assign T573 = T130[9:0];
  assign T130 = T131;
  assign T131 = {1'h0, Chain_1_io_ys_1};
  assign T574 = T132[9:0];
  assign T132 = T133;
  assign T133 = {1'h0, Chain_1_io_ys_2};
  assign T575 = T134[9:0];
  assign T134 = T135;
  assign T135 = {1'h0, Chain_1_io_ys_3};
  assign T576 = T136[9:0];
  assign T136 = T137;
  assign T137 = {1'h0, Chain_1_io_ys_4};
  assign T577 = T138[9:0];
  assign T138 = T139;
  assign T139 = {1'h0, Chain_1_io_ys_5};
  assign T578 = T140[9:0];
  assign T140 = T141;
  assign T141 = {1'h0, Chain_1_io_ys_6};
  assign T579 = T142[9:0];
  assign T142 = T143;
  assign T143 = {1'h0, Chain_1_io_ys_7};
  assign T580 = T144[9:0];
  assign T144 = T145;
  assign T145 = {1'h0, Chain_1_io_ys_8};
  assign T581 = T146[9:0];
  assign T146 = T147;
  assign T147 = {1'h0, Chain_1_io_ys_9};
  assign T582 = T148[9:0];
  assign T148 = T149;
  assign T149 = {1'h0, Chain_1_io_ys_10};
  assign T583 = T150[9:0];
  assign T150 = T151;
  assign T151 = {1'h0, Chain_1_io_ys_11};
  assign T584 = T152[9:0];
  assign T152 = T153;
  assign T153 = {1'h0, Chain_1_io_ys_12};
  assign T585 = T154[9:0];
  assign T154 = T155;
  assign T155 = {1'h0, Chain_1_io_ys_13};
  assign T586 = T156[9:0];
  assign T156 = T157;
  assign T157 = {1'h0, Chain_1_io_ys_14};
  assign T587 = T158[9:0];
  assign T158 = T159;
  assign T159 = {1'h0, Chain_1_io_ys_15};
  assign T588 = T160[9:0];
  assign T160 = T161;
  assign T161 = {1'h0, Chain_1_io_ys_16};
  assign T589 = T162[9:0];
  assign T162 = T163;
  assign T163 = {1'h0, Chain_1_io_ys_17};
  assign T590 = T164[9:0];
  assign T164 = T165;
  assign T165 = {1'h0, Chain_1_io_ys_18};
  assign T591 = T166[9:0];
  assign T166 = T167;
  assign T167 = {1'h0, Chain_1_io_ys_19};
  assign T592 = T168[9:0];
  assign T168 = T169;
  assign T169 = {1'h0, Chain_1_io_ys_20};
  assign T593 = T170[9:0];
  assign T170 = T171;
  assign T171 = {1'h0, Chain_1_io_ys_21};
  assign T594 = T172[9:0];
  assign T172 = T173;
  assign T173 = {1'h0, Chain_1_io_ys_22};
  assign T595 = T174[9:0];
  assign T174 = T175;
  assign T175 = {1'h0, Chain_1_io_ys_23};
  assign T596 = T176[9:0];
  assign T176 = T177;
  assign T177 = {1'h0, Chain_1_io_ys_24};
  assign T597 = T178[9:0];
  assign T178 = T179;
  assign T179 = {1'h0, Chain_1_io_ys_25};
  assign T598 = T180[9:0];
  assign T180 = T181;
  assign T181 = {1'h0, Chain_1_io_ys_26};
  assign T599 = T182[9:0];
  assign T182 = T183;
  assign T183 = {1'h0, Chain_1_io_ys_27};
  assign T600 = T184[9:0];
  assign T184 = T185;
  assign T185 = {1'h0, Chain_1_io_ys_28};
  assign T601 = T186[9:0];
  assign T186 = T187;
  assign T187 = {1'h0, Chain_1_io_ys_29};
  assign T602 = T188[9:0];
  assign T188 = T189;
  assign T189 = {1'h0, Chain_1_io_ys_30};
  assign T603 = T190[9:0];
  assign T190 = T191;
  assign T191 = {1'h0, Chain_1_io_ys_31};
  assign T604 = T192[9:0];
  assign T192 = T193;
  assign T193 = {1'h0, Chain_io_ys_0};
  assign T605 = T194[9:0];
  assign T194 = T195;
  assign T195 = {1'h0, Chain_io_ys_1};
  assign T606 = T196[9:0];
  assign T196 = T197;
  assign T197 = {1'h0, Chain_io_ys_2};
  assign T607 = T198[9:0];
  assign T198 = T199;
  assign T199 = {1'h0, Chain_io_ys_3};
  assign T608 = T200[9:0];
  assign T200 = T201;
  assign T201 = {1'h0, Chain_io_ys_4};
  assign T609 = T202[9:0];
  assign T202 = T203;
  assign T203 = {1'h0, Chain_io_ys_5};
  assign T610 = T204[9:0];
  assign T204 = T205;
  assign T205 = {1'h0, Chain_io_ys_6};
  assign T611 = T206[9:0];
  assign T206 = T207;
  assign T207 = {1'h0, Chain_io_ys_7};
  assign T612 = T208[9:0];
  assign T208 = T209;
  assign T209 = {1'h0, Chain_io_ys_8};
  assign T613 = T210[9:0];
  assign T210 = T211;
  assign T211 = {1'h0, Chain_io_ys_9};
  assign T614 = T212[9:0];
  assign T212 = T213;
  assign T213 = {1'h0, Chain_io_ys_10};
  assign T615 = T214[9:0];
  assign T214 = T215;
  assign T215 = {1'h0, Chain_io_ys_11};
  assign T616 = T216[9:0];
  assign T216 = T217;
  assign T217 = {1'h0, Chain_io_ys_12};
  assign T617 = T218[9:0];
  assign T218 = T219;
  assign T219 = {1'h0, Chain_io_ys_13};
  assign T618 = T220[9:0];
  assign T220 = T221;
  assign T221 = {1'h0, Chain_io_ys_14};
  assign T619 = T222[9:0];
  assign T222 = T223;
  assign T223 = {1'h0, Chain_io_ys_15};
  assign T620 = T224[9:0];
  assign T224 = T225;
  assign T225 = {1'h0, Chain_io_ys_16};
  assign T621 = T226[9:0];
  assign T226 = T227;
  assign T227 = {1'h0, Chain_io_ys_17};
  assign T622 = T228[9:0];
  assign T228 = T229;
  assign T229 = {1'h0, Chain_io_ys_18};
  assign T623 = T230[9:0];
  assign T230 = T231;
  assign T231 = {1'h0, Chain_io_ys_19};
  assign T624 = T232[9:0];
  assign T232 = T233;
  assign T233 = {1'h0, Chain_io_ys_20};
  assign T625 = T234[9:0];
  assign T234 = T235;
  assign T235 = {1'h0, Chain_io_ys_21};
  assign T626 = T236[9:0];
  assign T236 = T237;
  assign T237 = {1'h0, Chain_io_ys_22};
  assign T627 = T238[9:0];
  assign T238 = T239;
  assign T239 = {1'h0, Chain_io_ys_23};
  assign T628 = T240[9:0];
  assign T240 = T241;
  assign T241 = {1'h0, Chain_io_ys_24};
  assign T629 = T242[9:0];
  assign T242 = T243;
  assign T243 = {1'h0, Chain_io_ys_25};
  assign T630 = T244[9:0];
  assign T244 = T245;
  assign T245 = {1'h0, Chain_io_ys_26};
  assign T631 = T246[9:0];
  assign T246 = T247;
  assign T247 = {1'h0, Chain_io_ys_27};
  assign T632 = T248[9:0];
  assign T248 = T249;
  assign T249 = {1'h0, Chain_io_ys_28};
  assign T633 = T250[9:0];
  assign T250 = T251;
  assign T251 = {1'h0, Chain_io_ys_29};
  assign T634 = T252[9:0];
  assign T252 = T253;
  assign T253 = {1'h0, Chain_io_ys_30};
  assign T635 = T254[9:0];
  assign T254 = T255;
  assign T255 = {1'h0, Chain_io_ys_31};
  assign io_done = control_io_done;
  assign io_xOutValid = control_io_valid;
  assign io_xOut_0 = T256;
  assign T256 = T318 ? T288 : T257;
  assign T257 = T287 ? T273 : T258;
  assign T258 = T272 ? T266 : T259;
  assign T259 = T265 ? T263 : T260;
  assign T260 = T261 ? Activation_io_out_1 : Activation_io_out_0;
  assign T261 = T262[0];
  assign T262 = control_io_selectX;
  assign T263 = T264 ? Activation_io_out_3 : Activation_io_out_2;
  assign T264 = T262[0];
  assign T265 = T262[1];
  assign T266 = T271 ? T269 : T267;
  assign T267 = T268 ? Activation_io_out_5 : Activation_io_out_4;
  assign T268 = T262[0];
  assign T269 = T270 ? Activation_io_out_7 : Activation_io_out_6;
  assign T270 = T262[0];
  assign T271 = T262[1];
  assign T272 = T262[2];
  assign T273 = T286 ? T280 : T274;
  assign T274 = T279 ? T277 : T275;
  assign T275 = T276 ? Activation_io_out_9 : Activation_io_out_8;
  assign T276 = T262[0];
  assign T277 = T278 ? Activation_io_out_11 : Activation_io_out_10;
  assign T278 = T262[0];
  assign T279 = T262[1];
  assign T280 = T285 ? T283 : T281;
  assign T281 = T282 ? Activation_io_out_13 : Activation_io_out_12;
  assign T282 = T262[0];
  assign T283 = T284 ? Activation_io_out_15 : Activation_io_out_14;
  assign T284 = T262[0];
  assign T285 = T262[1];
  assign T286 = T262[2];
  assign T287 = T262[3];
  assign T288 = T317 ? T303 : T289;
  assign T289 = T302 ? T296 : T290;
  assign T290 = T295 ? T293 : T291;
  assign T291 = T292 ? Activation_io_out_17 : Activation_io_out_16;
  assign T292 = T262[0];
  assign T293 = T294 ? Activation_io_out_19 : Activation_io_out_18;
  assign T294 = T262[0];
  assign T295 = T262[1];
  assign T296 = T301 ? T299 : T297;
  assign T297 = T298 ? Activation_io_out_21 : Activation_io_out_20;
  assign T298 = T262[0];
  assign T299 = T300 ? Activation_io_out_23 : Activation_io_out_22;
  assign T300 = T262[0];
  assign T301 = T262[1];
  assign T302 = T262[2];
  assign T303 = T316 ? T310 : T304;
  assign T304 = T309 ? T307 : T305;
  assign T305 = T306 ? Activation_io_out_25 : Activation_io_out_24;
  assign T306 = T262[0];
  assign T307 = T308 ? Activation_io_out_27 : Activation_io_out_26;
  assign T308 = T262[0];
  assign T309 = T262[1];
  assign T310 = T315 ? T313 : T311;
  assign T311 = T312 ? Activation_io_out_29 : Activation_io_out_28;
  assign T312 = T262[0];
  assign T313 = T314 ? Activation_io_out_31 : Activation_io_out_30;
  assign T314 = T262[0];
  assign T315 = T262[1];
  assign T316 = T262[2];
  assign T317 = T262[3];
  assign T318 = T262[4];
  assign io_xOut_1 = T319;
  assign T319 = T381 ? T351 : T320;
  assign T320 = T350 ? T336 : T321;
  assign T321 = T335 ? T329 : T322;
  assign T322 = T328 ? T326 : T323;
  assign T323 = T324 ? Activation_1_io_out_1 : Activation_1_io_out_0;
  assign T324 = T325[0];
  assign T325 = control_io_selectX;
  assign T326 = T327 ? Activation_1_io_out_3 : Activation_1_io_out_2;
  assign T327 = T325[0];
  assign T328 = T325[1];
  assign T329 = T334 ? T332 : T330;
  assign T330 = T331 ? Activation_1_io_out_5 : Activation_1_io_out_4;
  assign T331 = T325[0];
  assign T332 = T333 ? Activation_1_io_out_7 : Activation_1_io_out_6;
  assign T333 = T325[0];
  assign T334 = T325[1];
  assign T335 = T325[2];
  assign T336 = T349 ? T343 : T337;
  assign T337 = T342 ? T340 : T338;
  assign T338 = T339 ? Activation_1_io_out_9 : Activation_1_io_out_8;
  assign T339 = T325[0];
  assign T340 = T341 ? Activation_1_io_out_11 : Activation_1_io_out_10;
  assign T341 = T325[0];
  assign T342 = T325[1];
  assign T343 = T348 ? T346 : T344;
  assign T344 = T345 ? Activation_1_io_out_13 : Activation_1_io_out_12;
  assign T345 = T325[0];
  assign T346 = T347 ? Activation_1_io_out_15 : Activation_1_io_out_14;
  assign T347 = T325[0];
  assign T348 = T325[1];
  assign T349 = T325[2];
  assign T350 = T325[3];
  assign T351 = T380 ? T366 : T352;
  assign T352 = T365 ? T359 : T353;
  assign T353 = T358 ? T356 : T354;
  assign T354 = T355 ? Activation_1_io_out_17 : Activation_1_io_out_16;
  assign T355 = T325[0];
  assign T356 = T357 ? Activation_1_io_out_19 : Activation_1_io_out_18;
  assign T357 = T325[0];
  assign T358 = T325[1];
  assign T359 = T364 ? T362 : T360;
  assign T360 = T361 ? Activation_1_io_out_21 : Activation_1_io_out_20;
  assign T361 = T325[0];
  assign T362 = T363 ? Activation_1_io_out_23 : Activation_1_io_out_22;
  assign T363 = T325[0];
  assign T364 = T325[1];
  assign T365 = T325[2];
  assign T366 = T379 ? T373 : T367;
  assign T367 = T372 ? T370 : T368;
  assign T368 = T369 ? Activation_1_io_out_25 : Activation_1_io_out_24;
  assign T369 = T325[0];
  assign T370 = T371 ? Activation_1_io_out_27 : Activation_1_io_out_26;
  assign T371 = T325[0];
  assign T372 = T325[1];
  assign T373 = T378 ? T376 : T374;
  assign T374 = T375 ? Activation_1_io_out_29 : Activation_1_io_out_28;
  assign T375 = T325[0];
  assign T376 = T377 ? Activation_1_io_out_31 : Activation_1_io_out_30;
  assign T377 = T325[0];
  assign T378 = T325[1];
  assign T379 = T325[2];
  assign T380 = T325[3];
  assign T381 = T325[4];
  assign io_xOut_2 = T382;
  assign T382 = T444 ? T414 : T383;
  assign T383 = T413 ? T399 : T384;
  assign T384 = T398 ? T392 : T385;
  assign T385 = T391 ? T389 : T386;
  assign T386 = T387 ? Activation_2_io_out_1 : Activation_2_io_out_0;
  assign T387 = T388[0];
  assign T388 = control_io_selectX;
  assign T389 = T390 ? Activation_2_io_out_3 : Activation_2_io_out_2;
  assign T390 = T388[0];
  assign T391 = T388[1];
  assign T392 = T397 ? T395 : T393;
  assign T393 = T394 ? Activation_2_io_out_5 : Activation_2_io_out_4;
  assign T394 = T388[0];
  assign T395 = T396 ? Activation_2_io_out_7 : Activation_2_io_out_6;
  assign T396 = T388[0];
  assign T397 = T388[1];
  assign T398 = T388[2];
  assign T399 = T412 ? T406 : T400;
  assign T400 = T405 ? T403 : T401;
  assign T401 = T402 ? Activation_2_io_out_9 : Activation_2_io_out_8;
  assign T402 = T388[0];
  assign T403 = T404 ? Activation_2_io_out_11 : Activation_2_io_out_10;
  assign T404 = T388[0];
  assign T405 = T388[1];
  assign T406 = T411 ? T409 : T407;
  assign T407 = T408 ? Activation_2_io_out_13 : Activation_2_io_out_12;
  assign T408 = T388[0];
  assign T409 = T410 ? Activation_2_io_out_15 : Activation_2_io_out_14;
  assign T410 = T388[0];
  assign T411 = T388[1];
  assign T412 = T388[2];
  assign T413 = T388[3];
  assign T414 = T443 ? T429 : T415;
  assign T415 = T428 ? T422 : T416;
  assign T416 = T421 ? T419 : T417;
  assign T417 = T418 ? Activation_2_io_out_17 : Activation_2_io_out_16;
  assign T418 = T388[0];
  assign T419 = T420 ? Activation_2_io_out_19 : Activation_2_io_out_18;
  assign T420 = T388[0];
  assign T421 = T388[1];
  assign T422 = T427 ? T425 : T423;
  assign T423 = T424 ? Activation_2_io_out_21 : Activation_2_io_out_20;
  assign T424 = T388[0];
  assign T425 = T426 ? Activation_2_io_out_23 : Activation_2_io_out_22;
  assign T426 = T388[0];
  assign T427 = T388[1];
  assign T428 = T388[2];
  assign T429 = T442 ? T436 : T430;
  assign T430 = T435 ? T433 : T431;
  assign T431 = T432 ? Activation_2_io_out_25 : Activation_2_io_out_24;
  assign T432 = T388[0];
  assign T433 = T434 ? Activation_2_io_out_27 : Activation_2_io_out_26;
  assign T434 = T388[0];
  assign T435 = T388[1];
  assign T436 = T441 ? T439 : T437;
  assign T437 = T438 ? Activation_2_io_out_29 : Activation_2_io_out_28;
  assign T438 = T388[0];
  assign T439 = T440 ? Activation_2_io_out_31 : Activation_2_io_out_30;
  assign T440 = T388[0];
  assign T441 = T388[1];
  assign T442 = T388[2];
  assign T443 = T388[3];
  assign T444 = T388[4];
  assign io_xOut_3 = T445;
  assign T445 = T507 ? T477 : T446;
  assign T446 = T476 ? T462 : T447;
  assign T447 = T461 ? T455 : T448;
  assign T448 = T454 ? T452 : T449;
  assign T449 = T450 ? Activation_3_io_out_1 : Activation_3_io_out_0;
  assign T450 = T451[0];
  assign T451 = control_io_selectX;
  assign T452 = T453 ? Activation_3_io_out_3 : Activation_3_io_out_2;
  assign T453 = T451[0];
  assign T454 = T451[1];
  assign T455 = T460 ? T458 : T456;
  assign T456 = T457 ? Activation_3_io_out_5 : Activation_3_io_out_4;
  assign T457 = T451[0];
  assign T458 = T459 ? Activation_3_io_out_7 : Activation_3_io_out_6;
  assign T459 = T451[0];
  assign T460 = T451[1];
  assign T461 = T451[2];
  assign T462 = T475 ? T469 : T463;
  assign T463 = T468 ? T466 : T464;
  assign T464 = T465 ? Activation_3_io_out_9 : Activation_3_io_out_8;
  assign T465 = T451[0];
  assign T466 = T467 ? Activation_3_io_out_11 : Activation_3_io_out_10;
  assign T467 = T451[0];
  assign T468 = T451[1];
  assign T469 = T474 ? T472 : T470;
  assign T470 = T471 ? Activation_3_io_out_13 : Activation_3_io_out_12;
  assign T471 = T451[0];
  assign T472 = T473 ? Activation_3_io_out_15 : Activation_3_io_out_14;
  assign T473 = T451[0];
  assign T474 = T451[1];
  assign T475 = T451[2];
  assign T476 = T451[3];
  assign T477 = T506 ? T492 : T478;
  assign T478 = T491 ? T485 : T479;
  assign T479 = T484 ? T482 : T480;
  assign T480 = T481 ? Activation_3_io_out_17 : Activation_3_io_out_16;
  assign T481 = T451[0];
  assign T482 = T483 ? Activation_3_io_out_19 : Activation_3_io_out_18;
  assign T483 = T451[0];
  assign T484 = T451[1];
  assign T485 = T490 ? T488 : T486;
  assign T486 = T487 ? Activation_3_io_out_21 : Activation_3_io_out_20;
  assign T487 = T451[0];
  assign T488 = T489 ? Activation_3_io_out_23 : Activation_3_io_out_22;
  assign T489 = T451[0];
  assign T490 = T451[1];
  assign T491 = T451[2];
  assign T492 = T505 ? T499 : T493;
  assign T493 = T498 ? T496 : T494;
  assign T494 = T495 ? Activation_3_io_out_25 : Activation_3_io_out_24;
  assign T495 = T451[0];
  assign T496 = T497 ? Activation_3_io_out_27 : Activation_3_io_out_26;
  assign T497 = T451[0];
  assign T498 = T451[1];
  assign T499 = T504 ? T502 : T500;
  assign T500 = T501 ? Activation_3_io_out_29 : Activation_3_io_out_28;
  assign T501 = T451[0];
  assign T502 = T503 ? Activation_3_io_out_31 : Activation_3_io_out_30;
  assign T503 = T451[0];
  assign T504 = T451[1];
  assign T505 = T451[2];
  assign T506 = T451[3];
  assign T507 = T451[4];
  assign io_startOut = io_start;
  assign io_ready = control_io_ready;
  WarpControl_0 control(.clk(clk), .reset(reset),
       .io_ready( control_io_ready ),
       .io_start( io_start ),
       .io_nextReady( io_pipeReady ),
       .io_valid( control_io_valid ),
       .io_done( control_io_done ),
       .io_selectX( control_io_selectX ),
       .io_memoryRestart( control_io_memoryRestart ),
       .io_chainRestart( control_io_chainRestart )
  );
  Chain_0 Chain(.clk(clk), .reset(reset),
       .io_weights_31( memoryStreamer_io_weights_31 ),
       .io_weights_30( memoryStreamer_io_weights_30 ),
       .io_weights_29( memoryStreamer_io_weights_29 ),
       .io_weights_28( memoryStreamer_io_weights_28 ),
       .io_weights_27( memoryStreamer_io_weights_27 ),
       .io_weights_26( memoryStreamer_io_weights_26 ),
       .io_weights_25( memoryStreamer_io_weights_25 ),
       .io_weights_24( memoryStreamer_io_weights_24 ),
       .io_weights_23( memoryStreamer_io_weights_23 ),
       .io_weights_22( memoryStreamer_io_weights_22 ),
       .io_weights_21( memoryStreamer_io_weights_21 ),
       .io_weights_20( memoryStreamer_io_weights_20 ),
       .io_weights_19( memoryStreamer_io_weights_19 ),
       .io_weights_18( memoryStreamer_io_weights_18 ),
       .io_weights_17( memoryStreamer_io_weights_17 ),
       .io_weights_16( memoryStreamer_io_weights_16 ),
       .io_weights_15( memoryStreamer_io_weights_15 ),
       .io_weights_14( memoryStreamer_io_weights_14 ),
       .io_weights_13( memoryStreamer_io_weights_13 ),
       .io_weights_12( memoryStreamer_io_weights_12 ),
       .io_weights_11( memoryStreamer_io_weights_11 ),
       .io_weights_10( memoryStreamer_io_weights_10 ),
       .io_weights_9( memoryStreamer_io_weights_9 ),
       .io_weights_8( memoryStreamer_io_weights_8 ),
       .io_weights_7( memoryStreamer_io_weights_7 ),
       .io_weights_6( memoryStreamer_io_weights_6 ),
       .io_weights_5( memoryStreamer_io_weights_5 ),
       .io_weights_4( memoryStreamer_io_weights_4 ),
       .io_weights_3( memoryStreamer_io_weights_3 ),
       .io_weights_2( memoryStreamer_io_weights_2 ),
       .io_weights_1( memoryStreamer_io_weights_1 ),
       .io_weights_0( memoryStreamer_io_weights_0 ),
       .io_bias( memoryStreamer_io_bias ),
       .io_restartIn( control_io_chainRestart ),
       .io_xs( io_xIn_0 ),
       .io_ys_31( Chain_io_ys_31 ),
       .io_ys_30( Chain_io_ys_30 ),
       .io_ys_29( Chain_io_ys_29 ),
       .io_ys_28( Chain_io_ys_28 ),
       .io_ys_27( Chain_io_ys_27 ),
       .io_ys_26( Chain_io_ys_26 ),
       .io_ys_25( Chain_io_ys_25 ),
       .io_ys_24( Chain_io_ys_24 ),
       .io_ys_23( Chain_io_ys_23 ),
       .io_ys_22( Chain_io_ys_22 ),
       .io_ys_21( Chain_io_ys_21 ),
       .io_ys_20( Chain_io_ys_20 ),
       .io_ys_19( Chain_io_ys_19 ),
       .io_ys_18( Chain_io_ys_18 ),
       .io_ys_17( Chain_io_ys_17 ),
       .io_ys_16( Chain_io_ys_16 ),
       .io_ys_15( Chain_io_ys_15 ),
       .io_ys_14( Chain_io_ys_14 ),
       .io_ys_13( Chain_io_ys_13 ),
       .io_ys_12( Chain_io_ys_12 ),
       .io_ys_11( Chain_io_ys_11 ),
       .io_ys_10( Chain_io_ys_10 ),
       .io_ys_9( Chain_io_ys_9 ),
       .io_ys_8( Chain_io_ys_8 ),
       .io_ys_7( Chain_io_ys_7 ),
       .io_ys_6( Chain_io_ys_6 ),
       .io_ys_5( Chain_io_ys_5 ),
       .io_ys_4( Chain_io_ys_4 ),
       .io_ys_3( Chain_io_ys_3 ),
       .io_ys_2( Chain_io_ys_2 ),
       .io_ys_1( Chain_io_ys_1 ),
       .io_ys_0( Chain_io_ys_0 )
  );
  Chain_0 Chain_1(.clk(clk), .reset(reset),
       .io_weights_31( memoryStreamer_io_weights_31 ),
       .io_weights_30( memoryStreamer_io_weights_30 ),
       .io_weights_29( memoryStreamer_io_weights_29 ),
       .io_weights_28( memoryStreamer_io_weights_28 ),
       .io_weights_27( memoryStreamer_io_weights_27 ),
       .io_weights_26( memoryStreamer_io_weights_26 ),
       .io_weights_25( memoryStreamer_io_weights_25 ),
       .io_weights_24( memoryStreamer_io_weights_24 ),
       .io_weights_23( memoryStreamer_io_weights_23 ),
       .io_weights_22( memoryStreamer_io_weights_22 ),
       .io_weights_21( memoryStreamer_io_weights_21 ),
       .io_weights_20( memoryStreamer_io_weights_20 ),
       .io_weights_19( memoryStreamer_io_weights_19 ),
       .io_weights_18( memoryStreamer_io_weights_18 ),
       .io_weights_17( memoryStreamer_io_weights_17 ),
       .io_weights_16( memoryStreamer_io_weights_16 ),
       .io_weights_15( memoryStreamer_io_weights_15 ),
       .io_weights_14( memoryStreamer_io_weights_14 ),
       .io_weights_13( memoryStreamer_io_weights_13 ),
       .io_weights_12( memoryStreamer_io_weights_12 ),
       .io_weights_11( memoryStreamer_io_weights_11 ),
       .io_weights_10( memoryStreamer_io_weights_10 ),
       .io_weights_9( memoryStreamer_io_weights_9 ),
       .io_weights_8( memoryStreamer_io_weights_8 ),
       .io_weights_7( memoryStreamer_io_weights_7 ),
       .io_weights_6( memoryStreamer_io_weights_6 ),
       .io_weights_5( memoryStreamer_io_weights_5 ),
       .io_weights_4( memoryStreamer_io_weights_4 ),
       .io_weights_3( memoryStreamer_io_weights_3 ),
       .io_weights_2( memoryStreamer_io_weights_2 ),
       .io_weights_1( memoryStreamer_io_weights_1 ),
       .io_weights_0( memoryStreamer_io_weights_0 ),
       .io_bias( memoryStreamer_io_bias ),
       .io_restartIn( control_io_chainRestart ),
       .io_xs( io_xIn_1 ),
       .io_ys_31( Chain_1_io_ys_31 ),
       .io_ys_30( Chain_1_io_ys_30 ),
       .io_ys_29( Chain_1_io_ys_29 ),
       .io_ys_28( Chain_1_io_ys_28 ),
       .io_ys_27( Chain_1_io_ys_27 ),
       .io_ys_26( Chain_1_io_ys_26 ),
       .io_ys_25( Chain_1_io_ys_25 ),
       .io_ys_24( Chain_1_io_ys_24 ),
       .io_ys_23( Chain_1_io_ys_23 ),
       .io_ys_22( Chain_1_io_ys_22 ),
       .io_ys_21( Chain_1_io_ys_21 ),
       .io_ys_20( Chain_1_io_ys_20 ),
       .io_ys_19( Chain_1_io_ys_19 ),
       .io_ys_18( Chain_1_io_ys_18 ),
       .io_ys_17( Chain_1_io_ys_17 ),
       .io_ys_16( Chain_1_io_ys_16 ),
       .io_ys_15( Chain_1_io_ys_15 ),
       .io_ys_14( Chain_1_io_ys_14 ),
       .io_ys_13( Chain_1_io_ys_13 ),
       .io_ys_12( Chain_1_io_ys_12 ),
       .io_ys_11( Chain_1_io_ys_11 ),
       .io_ys_10( Chain_1_io_ys_10 ),
       .io_ys_9( Chain_1_io_ys_9 ),
       .io_ys_8( Chain_1_io_ys_8 ),
       .io_ys_7( Chain_1_io_ys_7 ),
       .io_ys_6( Chain_1_io_ys_6 ),
       .io_ys_5( Chain_1_io_ys_5 ),
       .io_ys_4( Chain_1_io_ys_4 ),
       .io_ys_3( Chain_1_io_ys_3 ),
       .io_ys_2( Chain_1_io_ys_2 ),
       .io_ys_1( Chain_1_io_ys_1 ),
       .io_ys_0( Chain_1_io_ys_0 )
  );
  Chain_0 Chain_2(.clk(clk), .reset(reset),
       .io_weights_31( memoryStreamer_io_weights_31 ),
       .io_weights_30( memoryStreamer_io_weights_30 ),
       .io_weights_29( memoryStreamer_io_weights_29 ),
       .io_weights_28( memoryStreamer_io_weights_28 ),
       .io_weights_27( memoryStreamer_io_weights_27 ),
       .io_weights_26( memoryStreamer_io_weights_26 ),
       .io_weights_25( memoryStreamer_io_weights_25 ),
       .io_weights_24( memoryStreamer_io_weights_24 ),
       .io_weights_23( memoryStreamer_io_weights_23 ),
       .io_weights_22( memoryStreamer_io_weights_22 ),
       .io_weights_21( memoryStreamer_io_weights_21 ),
       .io_weights_20( memoryStreamer_io_weights_20 ),
       .io_weights_19( memoryStreamer_io_weights_19 ),
       .io_weights_18( memoryStreamer_io_weights_18 ),
       .io_weights_17( memoryStreamer_io_weights_17 ),
       .io_weights_16( memoryStreamer_io_weights_16 ),
       .io_weights_15( memoryStreamer_io_weights_15 ),
       .io_weights_14( memoryStreamer_io_weights_14 ),
       .io_weights_13( memoryStreamer_io_weights_13 ),
       .io_weights_12( memoryStreamer_io_weights_12 ),
       .io_weights_11( memoryStreamer_io_weights_11 ),
       .io_weights_10( memoryStreamer_io_weights_10 ),
       .io_weights_9( memoryStreamer_io_weights_9 ),
       .io_weights_8( memoryStreamer_io_weights_8 ),
       .io_weights_7( memoryStreamer_io_weights_7 ),
       .io_weights_6( memoryStreamer_io_weights_6 ),
       .io_weights_5( memoryStreamer_io_weights_5 ),
       .io_weights_4( memoryStreamer_io_weights_4 ),
       .io_weights_3( memoryStreamer_io_weights_3 ),
       .io_weights_2( memoryStreamer_io_weights_2 ),
       .io_weights_1( memoryStreamer_io_weights_1 ),
       .io_weights_0( memoryStreamer_io_weights_0 ),
       .io_bias( memoryStreamer_io_bias ),
       .io_restartIn( control_io_chainRestart ),
       .io_xs( io_xIn_2 ),
       .io_ys_31( Chain_2_io_ys_31 ),
       .io_ys_30( Chain_2_io_ys_30 ),
       .io_ys_29( Chain_2_io_ys_29 ),
       .io_ys_28( Chain_2_io_ys_28 ),
       .io_ys_27( Chain_2_io_ys_27 ),
       .io_ys_26( Chain_2_io_ys_26 ),
       .io_ys_25( Chain_2_io_ys_25 ),
       .io_ys_24( Chain_2_io_ys_24 ),
       .io_ys_23( Chain_2_io_ys_23 ),
       .io_ys_22( Chain_2_io_ys_22 ),
       .io_ys_21( Chain_2_io_ys_21 ),
       .io_ys_20( Chain_2_io_ys_20 ),
       .io_ys_19( Chain_2_io_ys_19 ),
       .io_ys_18( Chain_2_io_ys_18 ),
       .io_ys_17( Chain_2_io_ys_17 ),
       .io_ys_16( Chain_2_io_ys_16 ),
       .io_ys_15( Chain_2_io_ys_15 ),
       .io_ys_14( Chain_2_io_ys_14 ),
       .io_ys_13( Chain_2_io_ys_13 ),
       .io_ys_12( Chain_2_io_ys_12 ),
       .io_ys_11( Chain_2_io_ys_11 ),
       .io_ys_10( Chain_2_io_ys_10 ),
       .io_ys_9( Chain_2_io_ys_9 ),
       .io_ys_8( Chain_2_io_ys_8 ),
       .io_ys_7( Chain_2_io_ys_7 ),
       .io_ys_6( Chain_2_io_ys_6 ),
       .io_ys_5( Chain_2_io_ys_5 ),
       .io_ys_4( Chain_2_io_ys_4 ),
       .io_ys_3( Chain_2_io_ys_3 ),
       .io_ys_2( Chain_2_io_ys_2 ),
       .io_ys_1( Chain_2_io_ys_1 ),
       .io_ys_0( Chain_2_io_ys_0 )
  );
  Chain_0 Chain_3(.clk(clk), .reset(reset),
       .io_weights_31( memoryStreamer_io_weights_31 ),
       .io_weights_30( memoryStreamer_io_weights_30 ),
       .io_weights_29( memoryStreamer_io_weights_29 ),
       .io_weights_28( memoryStreamer_io_weights_28 ),
       .io_weights_27( memoryStreamer_io_weights_27 ),
       .io_weights_26( memoryStreamer_io_weights_26 ),
       .io_weights_25( memoryStreamer_io_weights_25 ),
       .io_weights_24( memoryStreamer_io_weights_24 ),
       .io_weights_23( memoryStreamer_io_weights_23 ),
       .io_weights_22( memoryStreamer_io_weights_22 ),
       .io_weights_21( memoryStreamer_io_weights_21 ),
       .io_weights_20( memoryStreamer_io_weights_20 ),
       .io_weights_19( memoryStreamer_io_weights_19 ),
       .io_weights_18( memoryStreamer_io_weights_18 ),
       .io_weights_17( memoryStreamer_io_weights_17 ),
       .io_weights_16( memoryStreamer_io_weights_16 ),
       .io_weights_15( memoryStreamer_io_weights_15 ),
       .io_weights_14( memoryStreamer_io_weights_14 ),
       .io_weights_13( memoryStreamer_io_weights_13 ),
       .io_weights_12( memoryStreamer_io_weights_12 ),
       .io_weights_11( memoryStreamer_io_weights_11 ),
       .io_weights_10( memoryStreamer_io_weights_10 ),
       .io_weights_9( memoryStreamer_io_weights_9 ),
       .io_weights_8( memoryStreamer_io_weights_8 ),
       .io_weights_7( memoryStreamer_io_weights_7 ),
       .io_weights_6( memoryStreamer_io_weights_6 ),
       .io_weights_5( memoryStreamer_io_weights_5 ),
       .io_weights_4( memoryStreamer_io_weights_4 ),
       .io_weights_3( memoryStreamer_io_weights_3 ),
       .io_weights_2( memoryStreamer_io_weights_2 ),
       .io_weights_1( memoryStreamer_io_weights_1 ),
       .io_weights_0( memoryStreamer_io_weights_0 ),
       .io_bias( memoryStreamer_io_bias ),
       .io_restartIn( control_io_chainRestart ),
       .io_xs( io_xIn_3 ),
       .io_ys_31( Chain_3_io_ys_31 ),
       .io_ys_30( Chain_3_io_ys_30 ),
       .io_ys_29( Chain_3_io_ys_29 ),
       .io_ys_28( Chain_3_io_ys_28 ),
       .io_ys_27( Chain_3_io_ys_27 ),
       .io_ys_26( Chain_3_io_ys_26 ),
       .io_ys_25( Chain_3_io_ys_25 ),
       .io_ys_24( Chain_3_io_ys_24 ),
       .io_ys_23( Chain_3_io_ys_23 ),
       .io_ys_22( Chain_3_io_ys_22 ),
       .io_ys_21( Chain_3_io_ys_21 ),
       .io_ys_20( Chain_3_io_ys_20 ),
       .io_ys_19( Chain_3_io_ys_19 ),
       .io_ys_18( Chain_3_io_ys_18 ),
       .io_ys_17( Chain_3_io_ys_17 ),
       .io_ys_16( Chain_3_io_ys_16 ),
       .io_ys_15( Chain_3_io_ys_15 ),
       .io_ys_14( Chain_3_io_ys_14 ),
       .io_ys_13( Chain_3_io_ys_13 ),
       .io_ys_12( Chain_3_io_ys_12 ),
       .io_ys_11( Chain_3_io_ys_11 ),
       .io_ys_10( Chain_3_io_ys_10 ),
       .io_ys_9( Chain_3_io_ys_9 ),
       .io_ys_8( Chain_3_io_ys_8 ),
       .io_ys_7( Chain_3_io_ys_7 ),
       .io_ys_6( Chain_3_io_ys_6 ),
       .io_ys_5( Chain_3_io_ys_5 ),
       .io_ys_4( Chain_3_io_ys_4 ),
       .io_ys_3( Chain_3_io_ys_3 ),
       .io_ys_2( Chain_3_io_ys_2 ),
       .io_ys_1( Chain_3_io_ys_1 ),
       .io_ys_0( Chain_3_io_ys_0 )
  );
  Activation_0 Activation(
       .io_in_31( T635 ),
       .io_in_30( T634 ),
       .io_in_29( T633 ),
       .io_in_28( T632 ),
       .io_in_27( T631 ),
       .io_in_26( T630 ),
       .io_in_25( T629 ),
       .io_in_24( T628 ),
       .io_in_23( T627 ),
       .io_in_22( T626 ),
       .io_in_21( T625 ),
       .io_in_20( T624 ),
       .io_in_19( T623 ),
       .io_in_18( T622 ),
       .io_in_17( T621 ),
       .io_in_16( T620 ),
       .io_in_15( T619 ),
       .io_in_14( T618 ),
       .io_in_13( T617 ),
       .io_in_12( T616 ),
       .io_in_11( T615 ),
       .io_in_10( T614 ),
       .io_in_9( T613 ),
       .io_in_8( T612 ),
       .io_in_7( T611 ),
       .io_in_6( T610 ),
       .io_in_5( T609 ),
       .io_in_4( T608 ),
       .io_in_3( T607 ),
       .io_in_2( T606 ),
       .io_in_1( T605 ),
       .io_in_0( T604 ),
       .io_out_31( Activation_io_out_31 ),
       .io_out_30( Activation_io_out_30 ),
       .io_out_29( Activation_io_out_29 ),
       .io_out_28( Activation_io_out_28 ),
       .io_out_27( Activation_io_out_27 ),
       .io_out_26( Activation_io_out_26 ),
       .io_out_25( Activation_io_out_25 ),
       .io_out_24( Activation_io_out_24 ),
       .io_out_23( Activation_io_out_23 ),
       .io_out_22( Activation_io_out_22 ),
       .io_out_21( Activation_io_out_21 ),
       .io_out_20( Activation_io_out_20 ),
       .io_out_19( Activation_io_out_19 ),
       .io_out_18( Activation_io_out_18 ),
       .io_out_17( Activation_io_out_17 ),
       .io_out_16( Activation_io_out_16 ),
       .io_out_15( Activation_io_out_15 ),
       .io_out_14( Activation_io_out_14 ),
       .io_out_13( Activation_io_out_13 ),
       .io_out_12( Activation_io_out_12 ),
       .io_out_11( Activation_io_out_11 ),
       .io_out_10( Activation_io_out_10 ),
       .io_out_9( Activation_io_out_9 ),
       .io_out_8( Activation_io_out_8 ),
       .io_out_7( Activation_io_out_7 ),
       .io_out_6( Activation_io_out_6 ),
       .io_out_5( Activation_io_out_5 ),
       .io_out_4( Activation_io_out_4 ),
       .io_out_3( Activation_io_out_3 ),
       .io_out_2( Activation_io_out_2 ),
       .io_out_1( Activation_io_out_1 ),
       .io_out_0( Activation_io_out_0 )
  );
  Activation_0 Activation_1(
       .io_in_31( T603 ),
       .io_in_30( T602 ),
       .io_in_29( T601 ),
       .io_in_28( T600 ),
       .io_in_27( T599 ),
       .io_in_26( T598 ),
       .io_in_25( T597 ),
       .io_in_24( T596 ),
       .io_in_23( T595 ),
       .io_in_22( T594 ),
       .io_in_21( T593 ),
       .io_in_20( T592 ),
       .io_in_19( T591 ),
       .io_in_18( T590 ),
       .io_in_17( T589 ),
       .io_in_16( T588 ),
       .io_in_15( T587 ),
       .io_in_14( T586 ),
       .io_in_13( T585 ),
       .io_in_12( T584 ),
       .io_in_11( T583 ),
       .io_in_10( T582 ),
       .io_in_9( T581 ),
       .io_in_8( T580 ),
       .io_in_7( T579 ),
       .io_in_6( T578 ),
       .io_in_5( T577 ),
       .io_in_4( T576 ),
       .io_in_3( T575 ),
       .io_in_2( T574 ),
       .io_in_1( T573 ),
       .io_in_0( T572 ),
       .io_out_31( Activation_1_io_out_31 ),
       .io_out_30( Activation_1_io_out_30 ),
       .io_out_29( Activation_1_io_out_29 ),
       .io_out_28( Activation_1_io_out_28 ),
       .io_out_27( Activation_1_io_out_27 ),
       .io_out_26( Activation_1_io_out_26 ),
       .io_out_25( Activation_1_io_out_25 ),
       .io_out_24( Activation_1_io_out_24 ),
       .io_out_23( Activation_1_io_out_23 ),
       .io_out_22( Activation_1_io_out_22 ),
       .io_out_21( Activation_1_io_out_21 ),
       .io_out_20( Activation_1_io_out_20 ),
       .io_out_19( Activation_1_io_out_19 ),
       .io_out_18( Activation_1_io_out_18 ),
       .io_out_17( Activation_1_io_out_17 ),
       .io_out_16( Activation_1_io_out_16 ),
       .io_out_15( Activation_1_io_out_15 ),
       .io_out_14( Activation_1_io_out_14 ),
       .io_out_13( Activation_1_io_out_13 ),
       .io_out_12( Activation_1_io_out_12 ),
       .io_out_11( Activation_1_io_out_11 ),
       .io_out_10( Activation_1_io_out_10 ),
       .io_out_9( Activation_1_io_out_9 ),
       .io_out_8( Activation_1_io_out_8 ),
       .io_out_7( Activation_1_io_out_7 ),
       .io_out_6( Activation_1_io_out_6 ),
       .io_out_5( Activation_1_io_out_5 ),
       .io_out_4( Activation_1_io_out_4 ),
       .io_out_3( Activation_1_io_out_3 ),
       .io_out_2( Activation_1_io_out_2 ),
       .io_out_1( Activation_1_io_out_1 ),
       .io_out_0( Activation_1_io_out_0 )
  );
  Activation_0 Activation_2(
       .io_in_31( T571 ),
       .io_in_30( T570 ),
       .io_in_29( T569 ),
       .io_in_28( T568 ),
       .io_in_27( T567 ),
       .io_in_26( T566 ),
       .io_in_25( T565 ),
       .io_in_24( T564 ),
       .io_in_23( T563 ),
       .io_in_22( T562 ),
       .io_in_21( T561 ),
       .io_in_20( T560 ),
       .io_in_19( T559 ),
       .io_in_18( T558 ),
       .io_in_17( T557 ),
       .io_in_16( T556 ),
       .io_in_15( T555 ),
       .io_in_14( T554 ),
       .io_in_13( T553 ),
       .io_in_12( T552 ),
       .io_in_11( T551 ),
       .io_in_10( T550 ),
       .io_in_9( T549 ),
       .io_in_8( T548 ),
       .io_in_7( T547 ),
       .io_in_6( T546 ),
       .io_in_5( T545 ),
       .io_in_4( T544 ),
       .io_in_3( T543 ),
       .io_in_2( T542 ),
       .io_in_1( T541 ),
       .io_in_0( T540 ),
       .io_out_31( Activation_2_io_out_31 ),
       .io_out_30( Activation_2_io_out_30 ),
       .io_out_29( Activation_2_io_out_29 ),
       .io_out_28( Activation_2_io_out_28 ),
       .io_out_27( Activation_2_io_out_27 ),
       .io_out_26( Activation_2_io_out_26 ),
       .io_out_25( Activation_2_io_out_25 ),
       .io_out_24( Activation_2_io_out_24 ),
       .io_out_23( Activation_2_io_out_23 ),
       .io_out_22( Activation_2_io_out_22 ),
       .io_out_21( Activation_2_io_out_21 ),
       .io_out_20( Activation_2_io_out_20 ),
       .io_out_19( Activation_2_io_out_19 ),
       .io_out_18( Activation_2_io_out_18 ),
       .io_out_17( Activation_2_io_out_17 ),
       .io_out_16( Activation_2_io_out_16 ),
       .io_out_15( Activation_2_io_out_15 ),
       .io_out_14( Activation_2_io_out_14 ),
       .io_out_13( Activation_2_io_out_13 ),
       .io_out_12( Activation_2_io_out_12 ),
       .io_out_11( Activation_2_io_out_11 ),
       .io_out_10( Activation_2_io_out_10 ),
       .io_out_9( Activation_2_io_out_9 ),
       .io_out_8( Activation_2_io_out_8 ),
       .io_out_7( Activation_2_io_out_7 ),
       .io_out_6( Activation_2_io_out_6 ),
       .io_out_5( Activation_2_io_out_5 ),
       .io_out_4( Activation_2_io_out_4 ),
       .io_out_3( Activation_2_io_out_3 ),
       .io_out_2( Activation_2_io_out_2 ),
       .io_out_1( Activation_2_io_out_1 ),
       .io_out_0( Activation_2_io_out_0 )
  );
  Activation_0 Activation_3(
       .io_in_31( T539 ),
       .io_in_30( T538 ),
       .io_in_29( T537 ),
       .io_in_28( T536 ),
       .io_in_27( T535 ),
       .io_in_26( T534 ),
       .io_in_25( T533 ),
       .io_in_24( T532 ),
       .io_in_23( T531 ),
       .io_in_22( T530 ),
       .io_in_21( T529 ),
       .io_in_20( T528 ),
       .io_in_19( T527 ),
       .io_in_18( T526 ),
       .io_in_17( T525 ),
       .io_in_16( T524 ),
       .io_in_15( T523 ),
       .io_in_14( T522 ),
       .io_in_13( T521 ),
       .io_in_12( T520 ),
       .io_in_11( T519 ),
       .io_in_10( T518 ),
       .io_in_9( T517 ),
       .io_in_8( T516 ),
       .io_in_7( T515 ),
       .io_in_6( T514 ),
       .io_in_5( T513 ),
       .io_in_4( T512 ),
       .io_in_3( T511 ),
       .io_in_2( T510 ),
       .io_in_1( T509 ),
       .io_in_0( T508 ),
       .io_out_31( Activation_3_io_out_31 ),
       .io_out_30( Activation_3_io_out_30 ),
       .io_out_29( Activation_3_io_out_29 ),
       .io_out_28( Activation_3_io_out_28 ),
       .io_out_27( Activation_3_io_out_27 ),
       .io_out_26( Activation_3_io_out_26 ),
       .io_out_25( Activation_3_io_out_25 ),
       .io_out_24( Activation_3_io_out_24 ),
       .io_out_23( Activation_3_io_out_23 ),
       .io_out_22( Activation_3_io_out_22 ),
       .io_out_21( Activation_3_io_out_21 ),
       .io_out_20( Activation_3_io_out_20 ),
       .io_out_19( Activation_3_io_out_19 ),
       .io_out_18( Activation_3_io_out_18 ),
       .io_out_17( Activation_3_io_out_17 ),
       .io_out_16( Activation_3_io_out_16 ),
       .io_out_15( Activation_3_io_out_15 ),
       .io_out_14( Activation_3_io_out_14 ),
       .io_out_13( Activation_3_io_out_13 ),
       .io_out_12( Activation_3_io_out_12 ),
       .io_out_11( Activation_3_io_out_11 ),
       .io_out_10( Activation_3_io_out_10 ),
       .io_out_9( Activation_3_io_out_9 ),
       .io_out_8( Activation_3_io_out_8 ),
       .io_out_7( Activation_3_io_out_7 ),
       .io_out_6( Activation_3_io_out_6 ),
       .io_out_5( Activation_3_io_out_5 ),
       .io_out_4( Activation_3_io_out_4 ),
       .io_out_3( Activation_3_io_out_3 ),
       .io_out_2( Activation_3_io_out_2 ),
       .io_out_1( Activation_3_io_out_1 ),
       .io_out_0( Activation_3_io_out_0 )
  );
  MemoryStreamer_0 memoryStreamer(.clk(clk), .reset(reset),
       .io_restart( control_io_memoryRestart ),
       .io_weights_31( memoryStreamer_io_weights_31 ),
       .io_weights_30( memoryStreamer_io_weights_30 ),
       .io_weights_29( memoryStreamer_io_weights_29 ),
       .io_weights_28( memoryStreamer_io_weights_28 ),
       .io_weights_27( memoryStreamer_io_weights_27 ),
       .io_weights_26( memoryStreamer_io_weights_26 ),
       .io_weights_25( memoryStreamer_io_weights_25 ),
       .io_weights_24( memoryStreamer_io_weights_24 ),
       .io_weights_23( memoryStreamer_io_weights_23 ),
       .io_weights_22( memoryStreamer_io_weights_22 ),
       .io_weights_21( memoryStreamer_io_weights_21 ),
       .io_weights_20( memoryStreamer_io_weights_20 ),
       .io_weights_19( memoryStreamer_io_weights_19 ),
       .io_weights_18( memoryStreamer_io_weights_18 ),
       .io_weights_17( memoryStreamer_io_weights_17 ),
       .io_weights_16( memoryStreamer_io_weights_16 ),
       .io_weights_15( memoryStreamer_io_weights_15 ),
       .io_weights_14( memoryStreamer_io_weights_14 ),
       .io_weights_13( memoryStreamer_io_weights_13 ),
       .io_weights_12( memoryStreamer_io_weights_12 ),
       .io_weights_11( memoryStreamer_io_weights_11 ),
       .io_weights_10( memoryStreamer_io_weights_10 ),
       .io_weights_9( memoryStreamer_io_weights_9 ),
       .io_weights_8( memoryStreamer_io_weights_8 ),
       .io_weights_7( memoryStreamer_io_weights_7 ),
       .io_weights_6( memoryStreamer_io_weights_6 ),
       .io_weights_5( memoryStreamer_io_weights_5 ),
       .io_weights_4( memoryStreamer_io_weights_4 ),
       .io_weights_3( memoryStreamer_io_weights_3 ),
       .io_weights_2( memoryStreamer_io_weights_2 ),
       .io_weights_1( memoryStreamer_io_weights_1 ),
       .io_weights_0( memoryStreamer_io_weights_0 ),
       .io_bias( memoryStreamer_io_bias )
  );
endmodule

module Counter_2(input clk, input reset,
    input  io_enable,
    input  io_rst,
    output[3:0] io_value
);

  reg [3:0] v;
  wire[3:0] T6;
  wire[3:0] T0;
  wire[3:0] T1;
  wire T2;
  wire[3:0] T3;
  wire T4;
  wire T5;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    v = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = v;
  assign T6 = reset ? 4'h0 : T0;
  assign T0 = T4 ? T3 : T1;
  assign T1 = T2 ? 4'h0 : v;
  assign T2 = io_enable & io_rst;
  assign T3 = v + 4'h1;
  assign T4 = io_enable & T5;
  assign T5 = io_rst ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      v <= 4'h0;
    end else if(T4) begin
      v <= T3;
    end else if(T2) begin
      v <= 4'h0;
    end
  end
endmodule

module Counter_5(input clk, input reset,
    input  io_enable,
    input  io_rst,
    output[7:0] io_value
);

  reg [7:0] v;
  wire[7:0] T6;
  wire[7:0] T0;
  wire[7:0] T1;
  wire T2;
  wire[7:0] T3;
  wire T4;
  wire T5;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    v = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = v;
  assign T6 = reset ? 8'h0 : T0;
  assign T0 = T4 ? T3 : T1;
  assign T1 = T2 ? 8'h0 : v;
  assign T2 = io_enable & io_rst;
  assign T3 = v + 8'h1;
  assign T4 = io_enable & T5;
  assign T5 = io_rst ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      v <= 8'h0;
    end else if(T4) begin
      v <= T3;
    end else if(T2) begin
      v <= 8'h0;
    end
  end
endmodule

module WarpControl_1(input clk, input reset,
    output io_ready,
    input  io_start,
    input  io_nextReady,
    output io_valid,
    output io_done,
    output[3:0] io_selectX,
    output io_memoryRestart,
    output io_chainRestart
);

  wire signalDone;
  reg  signalTailing;
  wire T8;
  wire signalLastActiveCycle;
  wire signalResetSelectX;
  reg  signalFirstOutputCycle;
  wire T9;
  wire signalOutputtingNext;
  wire T0;
  wire signalFirstReadyCycle;
  wire T1;
  wire signalLastCycleInPass;
  wire signalStartNewPass;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire[3:0] cycleInPass_io_value;
  wire[7:0] cycle_io_value;
  wire[3:0] tailCycle_io_value;
  wire[3:0] selectX_io_value;
  wire isActive_io_state;
  wire isReady_io_state;
  wire isOutputting_io_state;
  wire isTailing_io_state;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    signalTailing = {1{$random}};
    signalFirstOutputCycle = {1{$random}};
  end
// synthesis translate_on
`endif

  assign signalDone = tailCycle_io_value == 4'hf;
  assign T8 = reset ? 1'h0 : signalLastActiveCycle;
  assign signalLastActiveCycle = cycle_io_value == 8'hff;
  assign signalResetSelectX = selectX_io_value == 4'hf;
  assign T9 = reset ? 1'h0 : signalOutputtingNext;
  assign signalOutputtingNext = T0 & isActive_io_state;
  assign T0 = cycleInPass_io_value == 4'hf;
  assign signalFirstReadyCycle = T1 & isTailing_io_state;
  assign T1 = tailCycle_io_value == 4'h0;
  assign signalLastCycleInPass = cycleInPass_io_value == 4'hf;
  assign io_chainRestart = signalStartNewPass;
  assign signalStartNewPass = cycleInPass_io_value == 4'h0;
  assign io_memoryRestart = T2;
  assign T2 = T4 & T3;
  assign T3 = io_start ^ 1'h1;
  assign T4 = isReady_io_state | signalLastActiveCycle;
  assign io_selectX = selectX_io_value;
  assign io_done = signalDone;
  assign io_valid = isOutputting_io_state;
  assign io_ready = T5;
  assign T5 = T7 & T6;
  assign T6 = io_start ^ 1'h1;
  assign T7 = isReady_io_state & io_nextReady;
  Counter_2 cycleInPass(.clk(clk), .reset(reset),
       .io_enable( isActive_io_state ),
       .io_rst( signalLastCycleInPass ),
       .io_value( cycleInPass_io_value )
  );
  Counter_5 cycle(.clk(clk), .reset(reset),
       .io_enable( isActive_io_state ),
       .io_rst( signalLastActiveCycle ),
       .io_value( cycle_io_value )
  );
  Counter_2 tailCycle(.clk(clk), .reset(reset),
       .io_enable( isTailing_io_state ),
       .io_rst( signalDone ),
       .io_value( tailCycle_io_value )
  );
  Counter_2 selectX(.clk(clk), .reset(reset),
       .io_enable( isOutputting_io_state ),
       .io_rst( signalResetSelectX ),
       .io_value( selectX_io_value )
  );
  Switch_0 isActive(.clk(clk), .reset(reset),
       .io_signalOn( io_start ),
       .io_state( isActive_io_state ),
       .io_rst( signalLastActiveCycle )
  );
  Switch_1 isReady(.clk(clk), .reset(reset),
       .io_signalOn( signalFirstReadyCycle ),
       .io_state( isReady_io_state ),
       .io_rst( io_start )
  );
  Switch_0 isOutputting(.clk(clk), .reset(reset),
       .io_signalOn( signalFirstOutputCycle ),
       .io_state( isOutputting_io_state ),
       .io_rst( signalResetSelectX )
  );
  Switch_0 isTailing(.clk(clk), .reset(reset),
       .io_signalOn( signalTailing ),
       .io_state( isTailing_io_state ),
       .io_rst( signalDone )
  );

  always @(posedge clk) begin
    if(reset) begin
      signalTailing <= 1'h0;
    end else begin
      signalTailing <= signalLastActiveCycle;
    end
    if(reset) begin
      signalFirstOutputCycle <= 1'h0;
    end else begin
      signalFirstOutputCycle <= signalOutputtingNext;
    end
  end
endmodule

module Chain_1(input clk, input reset,
    input [15:0] io_weights_15,
    input [15:0] io_weights_14,
    input [15:0] io_weights_13,
    input [15:0] io_weights_12,
    input [15:0] io_weights_11,
    input [15:0] io_weights_10,
    input [15:0] io_weights_9,
    input [15:0] io_weights_8,
    input [15:0] io_weights_7,
    input [15:0] io_weights_6,
    input [15:0] io_weights_5,
    input [15:0] io_weights_4,
    input [15:0] io_weights_3,
    input [15:0] io_weights_2,
    input [15:0] io_weights_1,
    input [15:0] io_weights_0,
    input [7:0] io_bias,
    input  io_restartIn,
    input [15:0] io_xs,
    output[9:0] io_ys_15,
    output[9:0] io_ys_14,
    output[9:0] io_ys_13,
    output[9:0] io_ys_12,
    output[9:0] io_ys_11,
    output[9:0] io_ys_10,
    output[9:0] io_ys_9,
    output[9:0] io_ys_8,
    output[9:0] io_ys_7,
    output[9:0] io_ys_6,
    output[9:0] io_ys_5,
    output[9:0] io_ys_4,
    output[9:0] io_ys_3,
    output[9:0] io_ys_2,
    output[9:0] io_ys_1,
    output[9:0] io_ys_0
);

  wire[7:0] T32;
  wire[8:0] T0;
  wire[8:0] T1;
  wire[7:0] T33;
  wire[8:0] T2;
  wire[8:0] T3;
  wire[7:0] T34;
  wire[8:0] T4;
  wire[8:0] T5;
  wire[7:0] T35;
  wire[8:0] T6;
  wire[8:0] T7;
  wire[7:0] T36;
  wire[8:0] T8;
  wire[8:0] T9;
  wire[7:0] T37;
  wire[8:0] T10;
  wire[8:0] T11;
  wire[7:0] T38;
  wire[8:0] T12;
  wire[8:0] T13;
  wire[7:0] T39;
  wire[8:0] T14;
  wire[8:0] T15;
  wire[7:0] T40;
  wire[8:0] T16;
  wire[8:0] T17;
  wire[7:0] T41;
  wire[8:0] T18;
  wire[8:0] T19;
  wire[7:0] T42;
  wire[8:0] T20;
  wire[8:0] T21;
  wire[7:0] T43;
  wire[8:0] T22;
  wire[8:0] T23;
  wire[7:0] T44;
  wire[8:0] T24;
  wire[8:0] T25;
  wire[7:0] T45;
  wire[8:0] T26;
  wire[8:0] T27;
  wire[7:0] T46;
  wire[8:0] T28;
  wire[8:0] T29;
  wire[7:0] T47;
  wire[8:0] T30;
  wire[8:0] T31;
  wire[15:0] ProcessingUnit_io_xOut;
  wire[9:0] ProcessingUnit_io_yOut;
  wire ProcessingUnit_io_restartOut;
  wire[15:0] ProcessingUnit_1_io_xOut;
  wire[9:0] ProcessingUnit_1_io_yOut;
  wire ProcessingUnit_1_io_restartOut;
  wire[15:0] ProcessingUnit_2_io_xOut;
  wire[9:0] ProcessingUnit_2_io_yOut;
  wire ProcessingUnit_2_io_restartOut;
  wire[15:0] ProcessingUnit_3_io_xOut;
  wire[9:0] ProcessingUnit_3_io_yOut;
  wire ProcessingUnit_3_io_restartOut;
  wire[15:0] ProcessingUnit_4_io_xOut;
  wire[9:0] ProcessingUnit_4_io_yOut;
  wire ProcessingUnit_4_io_restartOut;
  wire[15:0] ProcessingUnit_5_io_xOut;
  wire[9:0] ProcessingUnit_5_io_yOut;
  wire ProcessingUnit_5_io_restartOut;
  wire[15:0] ProcessingUnit_6_io_xOut;
  wire[9:0] ProcessingUnit_6_io_yOut;
  wire ProcessingUnit_6_io_restartOut;
  wire[15:0] ProcessingUnit_7_io_xOut;
  wire[9:0] ProcessingUnit_7_io_yOut;
  wire ProcessingUnit_7_io_restartOut;
  wire[15:0] ProcessingUnit_8_io_xOut;
  wire[9:0] ProcessingUnit_8_io_yOut;
  wire ProcessingUnit_8_io_restartOut;
  wire[15:0] ProcessingUnit_9_io_xOut;
  wire[9:0] ProcessingUnit_9_io_yOut;
  wire ProcessingUnit_9_io_restartOut;
  wire[15:0] ProcessingUnit_10_io_xOut;
  wire[9:0] ProcessingUnit_10_io_yOut;
  wire ProcessingUnit_10_io_restartOut;
  wire[15:0] ProcessingUnit_11_io_xOut;
  wire[9:0] ProcessingUnit_11_io_yOut;
  wire ProcessingUnit_11_io_restartOut;
  wire[15:0] ProcessingUnit_12_io_xOut;
  wire[9:0] ProcessingUnit_12_io_yOut;
  wire ProcessingUnit_12_io_restartOut;
  wire[15:0] ProcessingUnit_13_io_xOut;
  wire[9:0] ProcessingUnit_13_io_yOut;
  wire ProcessingUnit_13_io_restartOut;
  wire[15:0] ProcessingUnit_14_io_xOut;
  wire[9:0] ProcessingUnit_14_io_yOut;
  wire ProcessingUnit_14_io_restartOut;
  wire[9:0] ProcessingUnit_15_io_yOut;


  assign T32 = T0[7:0];
  assign T0 = T1;
  assign T1 = {1'h0, io_bias};
  assign T33 = T2[7:0];
  assign T2 = T3;
  assign T3 = {1'h0, io_bias};
  assign T34 = T4[7:0];
  assign T4 = T5;
  assign T5 = {1'h0, io_bias};
  assign T35 = T6[7:0];
  assign T6 = T7;
  assign T7 = {1'h0, io_bias};
  assign T36 = T8[7:0];
  assign T8 = T9;
  assign T9 = {1'h0, io_bias};
  assign T37 = T10[7:0];
  assign T10 = T11;
  assign T11 = {1'h0, io_bias};
  assign T38 = T12[7:0];
  assign T12 = T13;
  assign T13 = {1'h0, io_bias};
  assign T39 = T14[7:0];
  assign T14 = T15;
  assign T15 = {1'h0, io_bias};
  assign T40 = T16[7:0];
  assign T16 = T17;
  assign T17 = {1'h0, io_bias};
  assign T41 = T18[7:0];
  assign T18 = T19;
  assign T19 = {1'h0, io_bias};
  assign T42 = T20[7:0];
  assign T20 = T21;
  assign T21 = {1'h0, io_bias};
  assign T43 = T22[7:0];
  assign T22 = T23;
  assign T23 = {1'h0, io_bias};
  assign T44 = T24[7:0];
  assign T24 = T25;
  assign T25 = {1'h0, io_bias};
  assign T45 = T26[7:0];
  assign T26 = T27;
  assign T27 = {1'h0, io_bias};
  assign T46 = T28[7:0];
  assign T28 = T29;
  assign T29 = {1'h0, io_bias};
  assign T47 = T30[7:0];
  assign T30 = T31;
  assign T31 = {1'h0, io_bias};
  assign io_ys_0 = ProcessingUnit_io_yOut;
  assign io_ys_1 = ProcessingUnit_1_io_yOut;
  assign io_ys_2 = ProcessingUnit_2_io_yOut;
  assign io_ys_3 = ProcessingUnit_3_io_yOut;
  assign io_ys_4 = ProcessingUnit_4_io_yOut;
  assign io_ys_5 = ProcessingUnit_5_io_yOut;
  assign io_ys_6 = ProcessingUnit_6_io_yOut;
  assign io_ys_7 = ProcessingUnit_7_io_yOut;
  assign io_ys_8 = ProcessingUnit_8_io_yOut;
  assign io_ys_9 = ProcessingUnit_9_io_yOut;
  assign io_ys_10 = ProcessingUnit_10_io_yOut;
  assign io_ys_11 = ProcessingUnit_11_io_yOut;
  assign io_ys_12 = ProcessingUnit_12_io_yOut;
  assign io_ys_13 = ProcessingUnit_13_io_yOut;
  assign io_ys_14 = ProcessingUnit_14_io_yOut;
  assign io_ys_15 = ProcessingUnit_15_io_yOut;
  ProcessingUnit ProcessingUnit(.clk(clk), .reset(reset),
       .io_xs( io_xs ),
       .io_ws( io_weights_0 ),
       .io_xOut( ProcessingUnit_io_xOut ),
       .io_yOut( ProcessingUnit_io_yOut ),
       .io_bias( T47 ),
       .io_restartIn( io_restartIn ),
       .io_restartOut( ProcessingUnit_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_1(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_io_xOut ),
       .io_ws( io_weights_1 ),
       .io_xOut( ProcessingUnit_1_io_xOut ),
       .io_yOut( ProcessingUnit_1_io_yOut ),
       .io_bias( T46 ),
       .io_restartIn( ProcessingUnit_io_restartOut ),
       .io_restartOut( ProcessingUnit_1_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_2(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_1_io_xOut ),
       .io_ws( io_weights_2 ),
       .io_xOut( ProcessingUnit_2_io_xOut ),
       .io_yOut( ProcessingUnit_2_io_yOut ),
       .io_bias( T45 ),
       .io_restartIn( ProcessingUnit_1_io_restartOut ),
       .io_restartOut( ProcessingUnit_2_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_3(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_2_io_xOut ),
       .io_ws( io_weights_3 ),
       .io_xOut( ProcessingUnit_3_io_xOut ),
       .io_yOut( ProcessingUnit_3_io_yOut ),
       .io_bias( T44 ),
       .io_restartIn( ProcessingUnit_2_io_restartOut ),
       .io_restartOut( ProcessingUnit_3_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_4(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_3_io_xOut ),
       .io_ws( io_weights_4 ),
       .io_xOut( ProcessingUnit_4_io_xOut ),
       .io_yOut( ProcessingUnit_4_io_yOut ),
       .io_bias( T43 ),
       .io_restartIn( ProcessingUnit_3_io_restartOut ),
       .io_restartOut( ProcessingUnit_4_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_5(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_4_io_xOut ),
       .io_ws( io_weights_5 ),
       .io_xOut( ProcessingUnit_5_io_xOut ),
       .io_yOut( ProcessingUnit_5_io_yOut ),
       .io_bias( T42 ),
       .io_restartIn( ProcessingUnit_4_io_restartOut ),
       .io_restartOut( ProcessingUnit_5_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_6(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_5_io_xOut ),
       .io_ws( io_weights_6 ),
       .io_xOut( ProcessingUnit_6_io_xOut ),
       .io_yOut( ProcessingUnit_6_io_yOut ),
       .io_bias( T41 ),
       .io_restartIn( ProcessingUnit_5_io_restartOut ),
       .io_restartOut( ProcessingUnit_6_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_7(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_6_io_xOut ),
       .io_ws( io_weights_7 ),
       .io_xOut( ProcessingUnit_7_io_xOut ),
       .io_yOut( ProcessingUnit_7_io_yOut ),
       .io_bias( T40 ),
       .io_restartIn( ProcessingUnit_6_io_restartOut ),
       .io_restartOut( ProcessingUnit_7_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_8(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_7_io_xOut ),
       .io_ws( io_weights_8 ),
       .io_xOut( ProcessingUnit_8_io_xOut ),
       .io_yOut( ProcessingUnit_8_io_yOut ),
       .io_bias( T39 ),
       .io_restartIn( ProcessingUnit_7_io_restartOut ),
       .io_restartOut( ProcessingUnit_8_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_9(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_8_io_xOut ),
       .io_ws( io_weights_9 ),
       .io_xOut( ProcessingUnit_9_io_xOut ),
       .io_yOut( ProcessingUnit_9_io_yOut ),
       .io_bias( T38 ),
       .io_restartIn( ProcessingUnit_8_io_restartOut ),
       .io_restartOut( ProcessingUnit_9_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_10(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_9_io_xOut ),
       .io_ws( io_weights_10 ),
       .io_xOut( ProcessingUnit_10_io_xOut ),
       .io_yOut( ProcessingUnit_10_io_yOut ),
       .io_bias( T37 ),
       .io_restartIn( ProcessingUnit_9_io_restartOut ),
       .io_restartOut( ProcessingUnit_10_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_11(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_10_io_xOut ),
       .io_ws( io_weights_11 ),
       .io_xOut( ProcessingUnit_11_io_xOut ),
       .io_yOut( ProcessingUnit_11_io_yOut ),
       .io_bias( T36 ),
       .io_restartIn( ProcessingUnit_10_io_restartOut ),
       .io_restartOut( ProcessingUnit_11_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_12(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_11_io_xOut ),
       .io_ws( io_weights_12 ),
       .io_xOut( ProcessingUnit_12_io_xOut ),
       .io_yOut( ProcessingUnit_12_io_yOut ),
       .io_bias( T35 ),
       .io_restartIn( ProcessingUnit_11_io_restartOut ),
       .io_restartOut( ProcessingUnit_12_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_13(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_12_io_xOut ),
       .io_ws( io_weights_13 ),
       .io_xOut( ProcessingUnit_13_io_xOut ),
       .io_yOut( ProcessingUnit_13_io_yOut ),
       .io_bias( T34 ),
       .io_restartIn( ProcessingUnit_12_io_restartOut ),
       .io_restartOut( ProcessingUnit_13_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_14(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_13_io_xOut ),
       .io_ws( io_weights_14 ),
       .io_xOut( ProcessingUnit_14_io_xOut ),
       .io_yOut( ProcessingUnit_14_io_yOut ),
       .io_bias( T33 ),
       .io_restartIn( ProcessingUnit_13_io_restartOut ),
       .io_restartOut( ProcessingUnit_14_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_15(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_14_io_xOut ),
       .io_ws( io_weights_15 ),
       //.io_xOut(  )
       .io_yOut( ProcessingUnit_15_io_yOut ),
       .io_bias( T32 ),
       .io_restartIn( ProcessingUnit_14_io_restartOut )
       //.io_restartOut(  )
  );
endmodule

module Activation_1(
    input [9:0] io_in_15,
    input [9:0] io_in_14,
    input [9:0] io_in_13,
    input [9:0] io_in_12,
    input [9:0] io_in_11,
    input [9:0] io_in_10,
    input [9:0] io_in_9,
    input [9:0] io_in_8,
    input [9:0] io_in_7,
    input [9:0] io_in_6,
    input [9:0] io_in_5,
    input [9:0] io_in_4,
    input [9:0] io_in_3,
    input [9:0] io_in_2,
    input [9:0] io_in_1,
    input [9:0] io_in_0,
    output io_out_15,
    output io_out_14,
    output io_out_13,
    output io_out_12,
    output io_out_11,
    output io_out_10,
    output io_out_9,
    output io_out_8,
    output io_out_7,
    output io_out_6,
    output io_out_5,
    output io_out_4,
    output io_out_3,
    output io_out_2,
    output io_out_1,
    output io_out_0
);

  wire T0;
  wire T1;
  wire[12:0] T2;
  wire[12:0] T3;
  wire T4;
  wire T5;
  wire[12:0] T6;
  wire[12:0] T7;
  wire T8;
  wire T9;
  wire[12:0] T10;
  wire[12:0] T11;
  wire T12;
  wire T13;
  wire[12:0] T14;
  wire[12:0] T15;
  wire T16;
  wire T17;
  wire[12:0] T18;
  wire[12:0] T19;
  wire T20;
  wire T21;
  wire[12:0] T22;
  wire[12:0] T23;
  wire T24;
  wire T25;
  wire[12:0] T26;
  wire[12:0] T27;
  wire T28;
  wire T29;
  wire[12:0] T30;
  wire[12:0] T31;
  wire T32;
  wire T33;
  wire[12:0] T34;
  wire[12:0] T35;
  wire T36;
  wire T37;
  wire[12:0] T38;
  wire[12:0] T39;
  wire T40;
  wire T41;
  wire[12:0] T42;
  wire[12:0] T43;
  wire T44;
  wire T45;
  wire[12:0] T46;
  wire[12:0] T47;
  wire T48;
  wire T49;
  wire[12:0] T50;
  wire[12:0] T51;
  wire T52;
  wire T53;
  wire[12:0] T54;
  wire[12:0] T55;
  wire T56;
  wire T57;
  wire[12:0] T58;
  wire[12:0] T59;
  wire T60;
  wire T61;
  wire[12:0] T62;
  wire[12:0] T63;


  assign io_out_0 = T0;
  assign T0 = ~ T1;
  assign T1 = T2[9];
  assign T2 = T3 - 13'h100;
  assign T3 = $signed(io_in_0) * $signed(3'h2);
  assign io_out_1 = T4;
  assign T4 = ~ T5;
  assign T5 = T6[9];
  assign T6 = T7 - 13'h100;
  assign T7 = $signed(io_in_1) * $signed(3'h2);
  assign io_out_2 = T8;
  assign T8 = ~ T9;
  assign T9 = T10[9];
  assign T10 = T11 - 13'h100;
  assign T11 = $signed(io_in_2) * $signed(3'h2);
  assign io_out_3 = T12;
  assign T12 = ~ T13;
  assign T13 = T14[9];
  assign T14 = T15 - 13'h100;
  assign T15 = $signed(io_in_3) * $signed(3'h2);
  assign io_out_4 = T16;
  assign T16 = ~ T17;
  assign T17 = T18[9];
  assign T18 = T19 - 13'h100;
  assign T19 = $signed(io_in_4) * $signed(3'h2);
  assign io_out_5 = T20;
  assign T20 = ~ T21;
  assign T21 = T22[9];
  assign T22 = T23 - 13'h100;
  assign T23 = $signed(io_in_5) * $signed(3'h2);
  assign io_out_6 = T24;
  assign T24 = ~ T25;
  assign T25 = T26[9];
  assign T26 = T27 - 13'h100;
  assign T27 = $signed(io_in_6) * $signed(3'h2);
  assign io_out_7 = T28;
  assign T28 = ~ T29;
  assign T29 = T30[9];
  assign T30 = T31 - 13'h100;
  assign T31 = $signed(io_in_7) * $signed(3'h2);
  assign io_out_8 = T32;
  assign T32 = ~ T33;
  assign T33 = T34[9];
  assign T34 = T35 - 13'h100;
  assign T35 = $signed(io_in_8) * $signed(3'h2);
  assign io_out_9 = T36;
  assign T36 = ~ T37;
  assign T37 = T38[9];
  assign T38 = T39 - 13'h100;
  assign T39 = $signed(io_in_9) * $signed(3'h2);
  assign io_out_10 = T40;
  assign T40 = ~ T41;
  assign T41 = T42[9];
  assign T42 = T43 - 13'h100;
  assign T43 = $signed(io_in_10) * $signed(3'h2);
  assign io_out_11 = T44;
  assign T44 = ~ T45;
  assign T45 = T46[9];
  assign T46 = T47 - 13'h100;
  assign T47 = $signed(io_in_11) * $signed(3'h2);
  assign io_out_12 = T48;
  assign T48 = ~ T49;
  assign T49 = T50[9];
  assign T50 = T51 - 13'h100;
  assign T51 = $signed(io_in_12) * $signed(3'h2);
  assign io_out_13 = T52;
  assign T52 = ~ T53;
  assign T53 = T54[9];
  assign T54 = T55 - 13'h100;
  assign T55 = $signed(io_in_13) * $signed(3'h2);
  assign io_out_14 = T56;
  assign T56 = ~ T57;
  assign T57 = T58[9];
  assign T58 = T59 - 13'h100;
  assign T59 = $signed(io_in_14) * $signed(3'h2);
  assign io_out_15 = T60;
  assign T60 = ~ T61;
  assign T61 = T62[9];
  assign T62 = T63 - 13'h100;
  assign T63 = $signed(io_in_15) * $signed(3'h2);
endmodule

module MemoryUnit_17(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[7:0] T5;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T6;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (T5)
    0: T0 = 32'h90d56b3d;
    1: T0 = 32'h3676111c;
    2: T0 = 32'heaff49bc;
    3: T0 = 32'h8602110e;
    4: T0 = 32'h28f73342;
    5: T0 = 32'hc63f3a9b;
    6: T0 = 32'h45b8f351;
    7: T0 = 32'hb0eb9c31;
    8: T0 = 32'h2126459;
    9: T0 = 32'h90e7f874;
    10: T0 = 32'hd92e80b8;
    11: T0 = 32'hcd541bee;
    12: T0 = 32'h553b0c81;
    13: T0 = 32'h663c8d96;
    14: T0 = 32'h4430b499;
    15: T0 = 32'h57263338;
    16: T0 = 32'h57a684fa;
    17: T0 = 32'h8d81e893;
    18: T0 = 32'h16cbdf8e;
    19: T0 = 32'h5098693b;
    20: T0 = 32'hb655c038;
    21: T0 = 32'hd9e8ebef;
    22: T0 = 32'hd334f13f;
    23: T0 = 32'hc6059a30;
    24: T0 = 32'hf1dc80d2;
    25: T0 = 32'heccfef7c;
    26: T0 = 32'h68b65916;
    27: T0 = 32'h27b5c0b;
    28: T0 = 32'hba3d627e;
    29: T0 = 32'hd969440a;
    30: T0 = 32'h6831f620;
    31: T0 = 32'h2bcbd9f4;
    32: T0 = 32'h3a5870dd;
    33: T0 = 32'h70b0979b;
    34: T0 = 32'h7d9f611;
    35: T0 = 32'h370ebe8a;
    36: T0 = 32'h5ac418c;
    37: T0 = 32'he54246d1;
    38: T0 = 32'h5a7f54ee;
    39: T0 = 32'h9cb03b4;
    40: T0 = 32'hcb949aaa;
    41: T0 = 32'h3623878f;
    42: T0 = 32'h1ddd12e;
    43: T0 = 32'hc4c07489;
    44: T0 = 32'h911157b7;
    45: T0 = 32'hdca57005;
    46: T0 = 32'he052ee66;
    47: T0 = 32'h8e85c8d5;
    48: T0 = 32'h8cd596aa;
    49: T0 = 32'hc6caace3;
    50: T0 = 32'h4fc37681;
    51: T0 = 32'h37dbfe88;
    52: T0 = 32'he556407f;
    53: T0 = 32'hddf20ad2;
    54: T0 = 32'h635019aa;
    55: T0 = 32'h8d8ac2d5;
    56: T0 = 32'h3a0ea272;
    57: T0 = 32'h9b158589;
    58: T0 = 32'h8db59de;
    59: T0 = 32'hbf70c8c9;
    60: T0 = 32'h4435c5f6;
    61: T0 = 32'hf5444437;
    62: T0 = 32'hf6e8afe7;
    63: T0 = 32'hb07d845;
    64: T0 = 32'h16dd22ac;
    65: T0 = 32'h10df3d8d;
    66: T0 = 32'h711ac911;
    67: T0 = 32'hfa6b544;
    68: T0 = 32'h69aa019f;
    69: T0 = 32'ha2113cc8;
    70: T0 = 32'h798fb2f6;
    71: T0 = 32'h6719c5f7;
    72: T0 = 32'hdf326761;
    73: T0 = 32'h2390b124;
    74: T0 = 32'h8b7ac4bc;
    75: T0 = 32'hd56c1fea;
    76: T0 = 32'hf3034a98;
    77: T0 = 32'h4510d76;
    78: T0 = 32'hc58ef49c;
    79: T0 = 32'hf685fa25;
    80: T0 = 32'hc93f7af6;
    81: T0 = 32'h5d47ed38;
    82: T0 = 32'hba34af65;
    83: T0 = 32'h8803298a;
    84: T0 = 32'h7a3b6300;
    85: T0 = 32'he295a4c8;
    86: T0 = 32'ha490b9be;
    87: T0 = 32'hc6141e23;
    88: T0 = 32'h6cb63252;
    89: T0 = 32'h4168876d;
    90: T0 = 32'hff22f534;
    91: T0 = 32'h56dfc583;
    92: T0 = 32'h27e126d7;
    93: T0 = 32'h225ad7cc;
    94: T0 = 32'h725ec94;
    95: T0 = 32'hf52e53ab;
    96: T0 = 32'h7b2ae626;
    97: T0 = 32'h5d5b80ec;
    98: T0 = 32'hef4262e1;
    99: T0 = 32'h916efd54;
    100: T0 = 32'h43e3283d;
    101: T0 = 32'hfec306da;
    102: T0 = 32'had25302e;
    103: T0 = 32'h27955724;
    104: T0 = 32'h1e5a8436;
    105: T0 = 32'h4b8d5d25;
    106: T0 = 32'h22d259b0;
    107: T0 = 32'hfe4549ca;
    108: T0 = 32'ha6665de7;
    109: T0 = 32'hf35804bc;
    110: T0 = 32'hbfe9b643;
    111: T0 = 32'h499c9796;
    112: T0 = 32'h670b80b8;
    113: T0 = 32'h12ce25cb;
    114: T0 = 32'h619e7bfd;
    115: T0 = 32'he7c49684;
    116: T0 = 32'h75bb9d6e;
    117: T0 = 32'h402c6b63;
    118: T0 = 32'he7ea11ea;
    119: T0 = 32'h30bf9308;
    120: T0 = 32'h9320b227;
    121: T0 = 32'ha8a201dd;
    122: T0 = 32'hbb3dfb03;
    123: T0 = 32'hdb26980a;
    124: T0 = 32'h588b9d79;
    125: T0 = 32'h363fa4db;
    126: T0 = 32'h44880741;
    127: T0 = 32'hb64785d5;
    128: T0 = 32'hc1b47a57;
    129: T0 = 32'h94e8a730;
    130: T0 = 32'heda33f25;
    131: T0 = 32'hf2815d8a;
    132: T0 = 32'hfe822504;
    133: T0 = 32'h41bfacc2;
    134: T0 = 32'hcbc01dbb;
    135: T0 = 32'h1da69f3b;
    136: T0 = 32'hf2c53fae;
    137: T0 = 32'h127203d9;
    138: T0 = 32'h8709fba2;
    139: T0 = 32'hf937e185;
    140: T0 = 32'hd44096c7;
    141: T0 = 32'h5574f3cc;
    142: T0 = 32'h57f8c05;
    143: T0 = 32'hfe7c449b;
    144: T0 = 32'hea474ce5;
    145: T0 = 32'hc8bbde22;
    146: T0 = 32'hb5c38603;
    147: T0 = 32'h7cbd78db;
    148: T0 = 32'hdec9ecf0;
    149: T0 = 32'h994847d1;
    150: T0 = 32'hcbe3cc6f;
    151: T0 = 32'h47bb5996;
    152: T0 = 32'hf1a482f8;
    153: T0 = 32'hb26a8fab;
    154: T0 = 32'h80dd445e;
    155: T0 = 32'h383b47b9;
    156: T0 = 32'ha81966fb;
    157: T0 = 32'h13eb6721;
    158: T0 = 32'hd9c1c626;
    159: T0 = 32'h2a6119ab;
    160: T0 = 32'h80511d1b;
    161: T0 = 32'h704fad5a;
    162: T0 = 32'he8b2804a;
    163: T0 = 32'hbf6247e1;
    164: T0 = 32'h68aafa73;
    165: T0 = 32'h6690ed27;
    166: T0 = 32'he4dc6f95;
    167: T0 = 32'h3dbbbe48;
    168: T0 = 32'h1b3acb8d;
    169: T0 = 32'h1ab022f2;
    170: T0 = 32'h13efbf4d;
    171: T0 = 32'hfd26c674;
    172: T0 = 32'hd5072a58;
    173: T0 = 32'ha6a7b669;
    174: T0 = 32'hd5e84b9c;
    175: T0 = 32'hc624668f;
    176: T0 = 32'h45bb37fe;
    177: T0 = 32'hc8812d99;
    178: T0 = 32'hd72afbfd;
    179: T0 = 32'h34965d12;
    180: T0 = 32'hf84b210c;
    181: T0 = 32'hd170b8c2;
    182: T0 = 32'h439239ba;
    183: T0 = 32'hcf0f9661;
    184: T0 = 32'h71a6e773;
    185: T0 = 32'hdb7aa77d;
    186: T0 = 32'h2c9679af;
    187: T0 = 32'h3478c8ce;
    188: T0 = 32'ha2b10afe;
    189: T0 = 32'h144b908e;
    190: T0 = 32'h7b25ecd1;
    191: T0 = 32'haa25e1ed;
    192: T0 = 32'h353978c7;
    193: T0 = 32'h76feb730;
    194: T0 = 32'h6b9cb402;
    195: T0 = 32'hab613eaa;
    196: T0 = 32'h5d8ae514;
    197: T0 = 32'h26050690;
    198: T0 = 32'h3cc9489e;
    199: T0 = 32'hb9dae99f;
    200: T0 = 32'h4e371b38;
    201: T0 = 32'h12b007cb;
    202: T0 = 32'h977fe5c6;
    203: T0 = 32'hed80a791;
    204: T0 = 32'h55429683;
    205: T0 = 32'h2694f347;
    206: T0 = 32'h95ceac2c;
    207: T0 = 32'h9c341c7b;
    208: T0 = 32'hcecf165e;
    209: T0 = 32'h846a7d9c;
    210: T0 = 32'h70cb8f6e;
    211: T0 = 32'h15fe412e;
    212: T0 = 32'h6179a20a;
    213: T0 = 32'hd86af98d;
    214: T0 = 32'h4bbff539;
    215: T0 = 32'hf4f99732;
    216: T0 = 32'h8b0a8895;
    217: T0 = 32'h88dfdb7c;
    218: T0 = 32'hc8b6cd46;
    219: T0 = 32'h34f5d07;
    220: T0 = 32'h1d3f04f6;
    221: T0 = 32'h213dc48a;
    222: T0 = 32'he48ad686;
    223: T0 = 32'h9282c1a4;
    224: T0 = 32'hd9f45ddb;
    225: T0 = 32'h5fffff50;
    226: T0 = 32'had1099ea;
    227: T0 = 32'h3bcd43a3;
    228: T0 = 32'h4122fac1;
    229: T0 = 32'h2510bd27;
    230: T0 = 32'hacc3e691;
    231: T0 = 32'had11be58;
    232: T0 = 32'h9e6ae3cc;
    233: T0 = 32'h778cab52;
    234: T0 = 32'h27d3f54d;
    235: T0 = 32'hfba56676;
    236: T0 = 32'heee6f35a;
    237: T0 = 32'ha25a9f69;
    238: T0 = 32'h97cc59bc;
    239: T0 = 32'h2cb1628b;
    240: T0 = 32'h642b6b62;
    241: T0 = 32'ha2b0b668;
    242: T0 = 32'h5497040;
    243: T0 = 32'h73b875f0;
    244: T0 = 32'h5edfe70;
    245: T0 = 32'hc96b8304;
    246: T0 = 32'hdbaf591d;
    247: T0 = 32'hbf3774b;
    248: T0 = 32'he3d98516;
    249: T0 = 32'h36576c89;
    250: T0 = 32'h19576b3;
    251: T0 = 32'h81b0c9e4;
    252: T0 = 32'hda25c1c7;
    253: T0 = 32'hcda012b1;
    254: T0 = 32'he8da29c3;
    255: T0 = 32'habd5342a;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[7:0];
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T6 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_18(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[7:0] T5;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T6;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (T5)
    0: T0 = 32'hccc76246;
    1: T0 = 32'h90cab2ec;
    2: T0 = 32'hb023e6c0;
    3: T0 = 32'hf6026777;
    4: T0 = 32'h76e96eb5;
    5: T0 = 32'hc998065c;
    6: T0 = 32'h435c1036;
    7: T0 = 32'h4adf7729;
    8: T0 = 32'h73919826;
    9: T0 = 32'h8bc05b0d;
    10: T0 = 32'h878b53f0;
    11: T0 = 32'h25ac58d4;
    12: T0 = 32'hf691dff7;
    13: T0 = 32'hd113262d;
    14: T0 = 32'h547735cb;
    15: T0 = 32'h89ee2616;
    16: T0 = 32'h981f58ef;
    17: T0 = 32'h1d282533;
    18: T0 = 32'hf0a77ee4;
    19: T0 = 32'h860acdaa;
    20: T0 = 32'h70792784;
    21: T0 = 32'hcafaeec4;
    22: T0 = 32'he7181d8a;
    23: T0 = 32'hf23d4b28;
    24: T0 = 32'h1c9217ba;
    25: T0 = 32'hc0da03c9;
    26: T0 = 32'hfda6fb3e;
    27: T0 = 32'h575fe883;
    28: T0 = 32'h243b8687;
    29: T0 = 32'h637bd304;
    30: T0 = 32'h4426ee65;
    31: T0 = 32'hc2b2045f;
    32: T0 = 32'hf3a23224;
    33: T0 = 32'h16fdb4a9;
    34: T0 = 32'h78b37480;
    35: T0 = 32'hc632b9a8;
    36: T0 = 32'hf939407a;
    37: T0 = 32'h5a2a0a9c;
    38: T0 = 32'hb9c55b7b;
    39: T0 = 32'hf63d5791;
    40: T0 = 32'hd232a6f2;
    41: T0 = 32'hc0f1cc8d;
    42: T0 = 32'hed6650ba;
    43: T0 = 32'h411f9989;
    44: T0 = 32'h747bc5a9;
    45: T0 = 32'h423e40b6;
    46: T0 = 32'h4430a6c3;
    47: T0 = 32'h76769b75;
    48: T0 = 32'hf9e47f47;
    49: T0 = 32'h3d749a34;
    50: T0 = 32'hda948618;
    51: T0 = 32'h113e687b;
    52: T0 = 32'h29ae72f1;
    53: T0 = 32'h967a34bc;
    54: T0 = 32'hb09dd414;
    55: T0 = 32'hb3d90c57;
    56: T0 = 32'h8c9b49d8;
    57: T0 = 32'h21d5fe0a;
    58: T0 = 32'h56f60488;
    59: T0 = 32'ha4325f2;
    60: T0 = 32'h992e6682;
    61: T0 = 32'h903b24;
    62: T0 = 32'hc5cafd3e;
    63: T0 = 32'hc2327b2a;
    64: T0 = 32'h95a92376;
    65: T0 = 32'h7c5e2f7c;
    66: T0 = 32'hf192a042;
    67: T0 = 32'h372426f4;
    68: T0 = 32'h69aa6677;
    69: T0 = 32'h6210142c;
    70: T0 = 32'hec8d31c0;
    71: T0 = 32'h753b0e5f;
    72: T0 = 32'h1b2a1f15;
    73: T0 = 32'h8907522;
    74: T0 = 32'hbfc4fc4;
    75: T0 = 32'he5265756;
    76: T0 = 32'hd5034c90;
    77: T0 = 32'h24f7af71;
    78: T0 = 32'hc1881d1f;
    79: T0 = 32'hee056f0f;
    80: T0 = 32'h51bfa2b6;
    81: T0 = 32'h104e35cb;
    82: T0 = 32'h209f79bc;
    83: T0 = 32'hcfe485ed;
    84: T0 = 32'h6dbf896a;
    85: T0 = 32'he2885b2f;
    86: T0 = 32'ha3ef1bfb;
    87: T0 = 32'h30bbc371;
    88: T0 = 32'h9720b6d7;
    89: T0 = 32'h88a2c0d5;
    90: T0 = 32'hdb7c83b2;
    91: T0 = 32'hc3269a4f;
    92: T0 = 32'h598b9da4;
    93: T0 = 32'h5637e0da;
    94: T0 = 32'hc48a0ac5;
    95: T0 = 32'hf6c780d5;
    96: T0 = 32'hc1b683a0;
    97: T0 = 32'h68860dc9;
    98: T0 = 32'hb77829bf;
    99: T0 = 32'h7c4697c4;
    100: T0 = 32'h26ef885b;
    101: T0 = 32'hf573193e;
    102: T0 = 32'hb3f1ae2;
    103: T0 = 32'h4bc1e0d5;
    104: T0 = 32'h6f9b7653;
    105: T0 = 32'h2b18b105;
    106: T0 = 32'hc2c4b8;
    107: T0 = 32'ha6e0db48;
    108: T0 = 32'hab956da0;
    109: T0 = 32'h9d810873;
    110: T0 = 32'h7b43adcd;
    111: T0 = 32'h9989b847;
    112: T0 = 32'h1c19bf5d;
    113: T0 = 32'hd749ca35;
    114: T0 = 32'hfaa4c011;
    115: T0 = 32'h8043fa53;
    116: T0 = 32'h695002b7;
    117: T0 = 32'h1abce4c8;
    118: T0 = 32'ha5b09c24;
    119: T0 = 32'hb63474c7;
    120: T0 = 32'h7e4258f8;
    121: T0 = 32'hc1f5fe62;
    122: T0 = 32'hfe201812;
    123: T0 = 32'h1d1f6f70;
    124: T0 = 32'h64ee60d6;
    125: T0 = 32'h627e2d3d;
    126: T0 = 32'h52cdc7e;
    127: T0 = 32'h53fafb2c;
    128: T0 = 32'hf322b4ed;
    129: T0 = 32'haf4c4bd3;
    130: T0 = 32'h854f691;
    131: T0 = 32'he9f1de83;
    132: T0 = 32'hc711011d;
    133: T0 = 32'h1f854c63;
    134: T0 = 32'hb46809aa;
    135: T0 = 32'hbe06f0c5;
    136: T0 = 32'hdc47127b;
    137: T0 = 32'h74350709;
    138: T0 = 32'h7d41d917;
    139: T0 = 32'h7a9d4851;
    140: T0 = 32'h4b6657de;
    141: T0 = 32'h4ada0551;
    142: T0 = 32'h8ebc7f75;
    143: T0 = 32'h7ddce8c5;
    144: T0 = 32'he70e313a;
    145: T0 = 32'h7c436fce;
    146: T0 = 32'h26fe994e;
    147: T0 = 32'h966407a4;
    148: T0 = 32'h2eaaca8f;
    149: T0 = 32'he6b0df2f;
    150: T0 = 32'h4d0431d6;
    151: T0 = 32'h3d99aab0;
    152: T0 = 32'h2f1ae729;
    153: T0 = 32'h1d843164;
    154: T0 = 32'h130bc785;
    155: T0 = 32'h4f27945a;
    156: T0 = 32'hf90f6b38;
    157: T0 = 32'hbfb58552;
    158: T0 = 32'h6341d59c;
    159: T0 = 32'h347edd7;
    160: T0 = 32'h8c8f958f;
    161: T0 = 32'h57bf0f53;
    162: T0 = 32'h6fd678f5;
    163: T0 = 32'h830bff84;
    164: T0 = 32'h911210d;
    165: T0 = 32'hc3bdd642;
    166: T0 = 32'h75e90a82;
    167: T0 = 32'ha4f4e06d;
    168: T0 = 32'h8076372b;
    169: T0 = 32'h446b05d9;
    170: T0 = 32'hbd76fabb;
    171: T0 = 32'hcd4daac0;
    172: T0 = 32'h447a9fc2;
    173: T0 = 32'h62349955;
    174: T0 = 32'h85222d6d;
    175: T0 = 32'h553cec4d;
    176: T0 = 32'heb86ef56;
    177: T0 = 32'h62a48a5c;
    178: T0 = 32'hb0ac097c;
    179: T0 = 32'h54804175;
    180: T0 = 32'hb87c3e62;
    181: T0 = 32'h40783127;
    182: T0 = 32'h2dc9711;
    183: T0 = 32'h5a7b3f4b;
    184: T0 = 32'h65323d8d;
    185: T0 = 32'ha4f25872;
    186: T0 = 32'hcda53fe3;
    187: T0 = 32'h40b85164;
    188: T0 = 32'h998bbdcb;
    189: T0 = 32'h8da5bb89;
    190: T0 = 32'h48160193;
    191: T0 = 32'h8ccb26a8;
    192: T0 = 32'h913432e6;
    193: T0 = 32'ha2a26f3e;
    194: T0 = 32'hdc32f24;
    195: T0 = 32'h319b1caa;
    196: T0 = 32'h87cd2607;
    197: T0 = 32'h8b5b34c9;
    198: T0 = 32'h192a3dde;
    199: T0 = 32'h1ae2ce33;
    200: T0 = 32'he2d523b3;
    201: T0 = 32'h36539549;
    202: T0 = 32'h9195cd70;
    203: T0 = 32'hc098ddca;
    204: T0 = 32'h984a86b4;
    205: T0 = 32'h7da4415e;
    206: T0 = 32'h88fbd41c;
    207: T0 = 32'hbdd5c9cf;
    208: T0 = 32'h9057a4b2;
    209: T0 = 32'h24511ecb;
    210: T0 = 32'hefe5016;
    211: T0 = 32'h866296ed;
    212: T0 = 32'h26ef99eb;
    213: T0 = 32'he6fb5b37;
    214: T0 = 32'h513d0be1;
    215: T0 = 32'h68d1e0d5;
    216: T0 = 32'h281b3643;
    217: T0 = 32'hb054085;
    218: T0 = 32'h520a8459;
    219: T0 = 32'hc6c59a18;
    220: T0 = 32'hd7179d18;
    221: T0 = 32'hec102973;
    222: T0 = 32'h6f611bcd;
    223: T0 = 32'h110e9c47;
    224: T0 = 32'he0f7ada;
    225: T0 = 32'h2625a358;
    226: T0 = 32'h52b5bbcc;
    227: T0 = 32'h4e3147a3;
    228: T0 = 32'hb81ab501;
    229: T0 = 32'h60bc6f27;
    230: T0 = 32'h1ad80989;
    231: T0 = 32'hd86abf6b;
    232: T0 = 32'h45b73e04;
    233: T0 = 32'h30f202db;
    234: T0 = 32'hcd0fbbe2;
    235: T0 = 32'h41bac264;
    236: T0 = 32'h3999bec7;
    237: T0 = 32'hc4a7b389;
    238: T0 = 32'h49360931;
    239: T0 = 32'he4e304db;
    240: T0 = 32'h9974fe73;
    241: T0 = 32'h36fe0a44;
    242: T0 = 32'h6fdcf27d;
    243: T0 = 32'heb64cf85;
    244: T0 = 32'h9d8abf35;
    245: T0 = 32'h261f8123;
    246: T0 = 32'h584b0d08;
    247: T0 = 32'h39ea3e4f;
    248: T0 = 32'h8a5f1d35;
    249: T0 = 32'h36375e59;
    250: T0 = 32'hd359ba17;
    251: T0 = 32'hed344954;
    252: T0 = 32'h59428d52;
    253: T0 = 32'hcb4b3c9;
    254: T0 = 32'h85c31971;
    255: T0 = 32'h9e35260f;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[7:0];
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T6 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_19(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[7:0] T5;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T6;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (T5)
    0: T0 = 32'h37387f55;
    1: T0 = 32'hee510b1c;
    2: T0 = 32'hde762b35;
    3: T0 = 32'h6134146;
    4: T0 = 32'h6ad72683;
    5: T0 = 32'hfefab097;
    6: T0 = 32'h51149519;
    7: T0 = 32'hcc0c946b;
    8: T0 = 32'h7a0f2d85;
    9: T0 = 32'h1b05737c;
    10: T0 = 32'h4e2b9fe1;
    11: T0 = 32'h3e48f156;
    12: T0 = 32'h67359ec6;
    13: T0 = 32'hf4c1bbc8;
    14: T0 = 32'h6bad0511;
    15: T0 = 32'h32e77a0;
    16: T0 = 32'h17075ced;
    17: T0 = 32'h1198f932;
    18: T0 = 32'h759bc613;
    19: T0 = 32'h9d0af8b9;
    20: T0 = 32'h76bc190;
    21: T0 = 32'hc18be6d5;
    22: T0 = 32'hffa7ce77;
    23: T0 = 32'he0d74896;
    24: T0 = 32'ha9b443f8;
    25: T0 = 32'hca49afaa;
    26: T0 = 32'ha1f4645a;
    27: T0 = 32'h846d2791;
    28: T0 = 32'ha63b6692;
    29: T0 = 32'h7a184924;
    30: T0 = 32'hec63e6ee;
    31: T0 = 32'hd68cbb2b;
    32: T0 = 32'hcbd1877a;
    33: T0 = 32'h324a68c7;
    34: T0 = 32'h609fc9c9;
    35: T0 = 32'hb7c4e191;
    36: T0 = 32'h7dabd83c;
    37: T0 = 32'h2208ed6d;
    38: T0 = 32'habeb36a1;
    39: T0 = 32'h31bb52e8;
    40: T0 = 32'hb320c4ee;
    41: T0 = 32'h88e2f8b4;
    42: T0 = 32'h9b7cdb1f;
    43: T0 = 32'h5106486e;
    44: T0 = 32'h588b7378;
    45: T0 = 32'h16378cb8;
    46: T0 = 32'h40887352;
    47: T0 = 32'hf6c7e3e6;
    48: T0 = 32'hc1b687db;
    49: T0 = 32'h300269cb;
    50: T0 = 32'ha75ed9fc;
    51: T0 = 32'haaecdeaf;
    52: T0 = 32'h6ae1d8a;
    53: T0 = 32'h6626eb63;
    54: T0 = 32'h4e2e3591;
    55: T0 = 32'h39cab028;
    56: T0 = 32'h8b1abf8f;
    57: T0 = 32'h3b052070;
    58: T0 = 32'h53d9bb07;
    59: T0 = 32'hefa4b84f;
    60: T0 = 32'hd916933e;
    61: T0 = 32'hbc35b6cb;
    62: T0 = 32'hb6c35751;
    63: T0 = 32'h1f11e5c5;
    64: T0 = 32'hccde16eb;
    65: T0 = 32'h5b28f8b3;
    66: T0 = 32'h3428cfb4;
    67: T0 = 32'h19aa593b;
    68: T0 = 32'h2134c0f8;
    69: T0 = 32'hf162e9c1;
    70: T0 = 32'hbb8cb63f;
    71: T0 = 32'heb519270;
    72: T0 = 32'h8771c0f2;
    73: T0 = 32'he7d5fd7d;
    74: T0 = 32'ha8d0591f;
    75: T0 = 32'h60e95cbb;
    76: T0 = 32'h87e6027e;
    77: T0 = 32'hc00944ae;
    78: T0 = 32'h98bef6e6;
    79: T0 = 32'ha89af1e4;
    80: T0 = 32'hb379fe5d;
    81: T0 = 32'hcb08ca16;
    82: T0 = 32'h11c90f9d;
    83: T0 = 32'h59bce81a;
    84: T0 = 32'h83256304;
    85: T0 = 32'h9dc864c3;
    86: T0 = 32'h9bbfb40a;
    87: T0 = 32'h5739d826;
    88: T0 = 32'h91a819b8;
    89: T0 = 32'hbe8bd77a;
    90: T0 = 32'h60b4f976;
    91: T0 = 32'h90a97743;
    92: T0 = 32'h882d42d6;
    93: T0 = 32'h9b69d7ac;
    94: T0 = 32'hf8defe71;
    95: T0 = 32'h23c15bf9;
    96: T0 = 32'hb15894aa;
    97: T0 = 32'h5d9bad33;
    98: T0 = 32'h7d50f2c1;
    99: T0 = 32'h998ebe88;
    100: T0 = 32'h43ab413d;
    101: T0 = 32'hb3c343c0;
    102: T0 = 32'hbd2329a6;
    103: T0 = 32'ha695e2c4;
    104: T0 = 32'haa59d27a;
    105: T0 = 32'h674c8f89;
    106: T0 = 32'hb3d0797f;
    107: T0 = 32'he40fc4c0;
    108: T0 = 32'ha676d574;
    109: T0 = 32'h63181077;
    110: T0 = 32'h9df8ac7c;
    111: T0 = 32'h59fccac7;
    112: T0 = 32'h6acbef5d;
    113: T0 = 32'h69070a1c;
    114: T0 = 32'h30ac69bd;
    115: T0 = 32'h19ee4954;
    116: T0 = 32'h217c3705;
    117: T0 = 32'hfee0b48b;
    118: T0 = 32'hb2bcfe04;
    119: T0 = 32'hf655557f;
    120: T0 = 32'hd3a7d15;
    121: T0 = 32'hed9d7c70;
    122: T0 = 32'h68f6bca0;
    123: T0 = 32'h26e973e6;
    124: T0 = 32'hb3ad0cc0;
    125: T0 = 32'haa29bb98;
    126: T0 = 32'hba807db9;
    127: T0 = 32'h19a76a4;
    128: T0 = 32'h26b88ba8;
    129: T0 = 32'h5a76c405;
    130: T0 = 32'hab1879bf;
    131: T0 = 32'hab68f155;
    132: T0 = 32'h45a29956;
    133: T0 = 32'h6615f0db;
    134: T0 = 32'h259bc22e;
    135: T0 = 32'h399851e5;
    136: T0 = 32'he2ae27b;
    137: T0 = 32'h2306a4b4;
    138: T0 = 32'h1b58b078;
    139: T0 = 32'hfdc4a6f8;
    140: T0 = 32'hc5c644cb;
    141: T0 = 32'h6ed668fe;
    142: T0 = 32'h97a8f0ba;
    143: T0 = 32'h369db330;
    144: T0 = 32'h67abcda1;
    145: T0 = 32'haf6d8e66;
    146: T0 = 32'hd825a003;
    147: T0 = 32'h40b13ed5;
    148: T0 = 32'hf951edf7;
    149: T0 = 32'h19784670;
    150: T0 = 32'ha0c00ac6;
    151: T0 = 32'hd72e60cf;
    152: T0 = 32'h7465536d;
    153: T0 = 32'ha0f07e83;
    154: T0 = 32'hfe2956dd;
    155: T0 = 32'h18ba27f8;
    156: T0 = 32'h6ee07158;
    157: T0 = 32'h4c22f35;
    158: T0 = 32'h29bd1d3e;
    159: T0 = 32'h60626e43;
    160: T0 = 32'h33205d47;
    161: T0 = 32'hb4fafa34;
    162: T0 = 32'h6edb8e03;
    163: T0 = 32'hd2647a3b;
    164: T0 = 32'h9eed6214;
    165: T0 = 32'hce5b24d0;
    166: T0 = 32'h496ff434;
    167: T0 = 32'h31f97c96;
    168: T0 = 32'haa1869f8;
    169: T0 = 32'h86f7ff2a;
    170: T0 = 32'hd53c76df;
    171: T0 = 32'hc73727e0;
    172: T0 = 32'hd91b729a;
    173: T0 = 32'h453c1725;
    174: T0 = 32'hc45371ae;
    175: T0 = 32'h13456b0a;
    176: T0 = 32'hc9c73d20;
    177: T0 = 32'ha6584d47;
    178: T0 = 32'h4a5699ab;
    179: T0 = 32'h336b1c4;
    180: T0 = 32'h8ecfc47a;
    181: T0 = 32'h8e6bffd8;
    182: T0 = 32'h5927b1ea;
    183: T0 = 32'ha5c0c8d6;
    184: T0 = 32'hea5f36db;
    185: T0 = 32'h92595f4;
    186: T0 = 32'h55724c33;
    187: T0 = 32'hcf428d6a;
    188: T0 = 32'h795e68bc;
    189: T0 = 32'hc108c7a;
    190: T0 = 32'ha553c6f2;
    191: T0 = 32'h517db0d3;
    192: T0 = 32'hcf8780aa;
    193: T0 = 32'h10a2f5e3;
    194: T0 = 32'ha7fbd642;
    195: T0 = 32'hb64266a9;
    196: T0 = 32'hb6a8c8b8;
    197: T0 = 32'he6b04774;
    198: T0 = 32'h47744cbf;
    199: T0 = 32'h39db2b98;
    200: T0 = 32'h4b9a93ea;
    201: T0 = 32'ha76a898b;
    202: T0 = 32'h818d6b1e;
    203: T0 = 32'h434f8409;
    204: T0 = 32'h840bf33f;
    205: T0 = 32'he73c5463;
    206: T0 = 32'hc663aa66;
    207: T0 = 32'h78688df;
    208: T0 = 32'hc9df337e;
    209: T0 = 32'ha1b00d9c;
    210: T0 = 32'h5cb6bfc;
    211: T0 = 32'h319b411e;
    212: T0 = 32'h87c4330c;
    213: T0 = 32'h8d7eb8cb;
    214: T0 = 32'h9befb138;
    215: T0 = 32'hbeb9721;
    216: T0 = 32'hc3cceed7;
    217: T0 = 32'hb607a378;
    218: T0 = 32'h195bba0;
    219: T0 = 32'hcaf1f8ee;
    220: T0 = 32'hda680cf7;
    221: T0 = 32'hdde5908a;
    222: T0 = 32'hacfba6d1;
    223: T0 = 32'hdd7e3a1;
    224: T0 = 32'ha4d76ad5;
    225: T0 = 32'h977cb738;
    226: T0 = 32'hc8963626;
    227: T0 = 32'h23bb1a0a;
    228: T0 = 32'hc91127a5;
    229: T0 = 32'ha0c34d3;
    230: T0 = 32'hf4c2cddc;
    231: T0 = 32'hb42e0927;
    232: T0 = 32'hd0657b18;
    233: T0 = 32'h50e706cb;
    234: T0 = 32'hff7cb7e0;
    235: T0 = 32'h5917e7b5;
    236: T0 = 32'h596eaec3;
    237: T0 = 32'h627ef347;
    238: T0 = 32'h84b8aeb4;
    239: T0 = 32'h67701c39;
    240: T0 = 32'hf3e47e75;
    241: T0 = 32'h49018f54;
    242: T0 = 32'hd025a861;
    243: T0 = 32'h549b298a;
    244: T0 = 32'h61542527;
    245: T0 = 32'hf9e074d3;
    246: T0 = 32'hb714ac62;
    247: T0 = 32'hc23d8c5f;
    248: T0 = 32'h3580363d;
    249: T0 = 32'hc8ce1756;
    250: T0 = 32'haca5eeb6;
    251: T0 = 32'h14ef4d76;
    252: T0 = 32'ha6ad6e94;
    253: T0 = 32'h734bbbe8;
    254: T0 = 32'h68ac9c31;
    255: T0 = 32'h3ca5eab;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[7:0];
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T6 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_20(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[7:0] T5;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T6;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (T5)
    0: T0 = 32'hc95558a6;
    1: T0 = 32'ha459070a;
    2: T0 = 32'h5a963702;
    3: T0 = 32'h413eb68c;
    4: T0 = 32'h8acfe156;
    5: T0 = 32'h9bcb5fda;
    6: T0 = 32'h596709ea;
    7: T0 = 32'hc401e995;
    8: T0 = 32'hf8573661;
    9: T0 = 32'h7c250599;
    10: T0 = 32'h4276e4d8;
    11: T0 = 32'h8c428291;
    12: T0 = 32'hff59dc85;
    13: T0 = 32'h1d00d077;
    14: T0 = 32'hedd9bd8d;
    15: T0 = 32'h53751c5b;
    16: T0 = 32'h44c4b4aa;
    17: T0 = 32'h3aa6ad63;
    18: T0 = 32'h2f7cf281;
    19: T0 = 32'ha240fc80;
    20: T0 = 32'h25ee487e;
    21: T0 = 32'he7f74048;
    22: T0 = 32'h143c09aa;
    23: T0 = 32'h29c0c2c5;
    24: T0 = 32'he1f9272;
    25: T0 = 32'h17558789;
    26: T0 = 32'h3d025098;
    27: T0 = 32'h4fd4c8c8;
    28: T0 = 32'h57c6c4c6;
    29: T0 = 32'h4c944077;
    30: T0 = 32'h25b0aeef;
    31: T0 = 32'h1d9e9847;
    32: T0 = 32'h1a2f6b05;
    33: T0 = 32'h85d91f6c;
    34: T0 = 32'h4f873875;
    35: T0 = 32'h97b7bfe5;
    36: T0 = 32'heecf3fe7;
    37: T0 = 32'hcd8d142c;
    38: T0 = 32'h67f34e40;
    39: T0 = 32'h448e45df;
    40: T0 = 32'ha8967f09;
    41: T0 = 32'h5a283000;
    42: T0 = 32'h3fa26a9;
    43: T0 = 32'h8d44a3e4;
    44: T0 = 32'h361b9d89;
    45: T0 = 32'hf33cbb75;
    46: T0 = 32'he57529d9;
    47: T0 = 32'h5a643e1b;
    48: T0 = 32'hcdc75d1b;
    49: T0 = 32'h84b87a32;
    50: T0 = 32'h4ab7894a;
    51: T0 = 32'h80db4339;
    52: T0 = 32'h685ffa81;
    53: T0 = 32'hd87bf525;
    54: T0 = 32'h517de614;
    55: T0 = 32'hc226287a;
    56: T0 = 32'h98c64bc8;
    57: T0 = 32'hc4f1b962;
    58: T0 = 32'hfc26644d;
    59: T0 = 32'h185c6666;
    60: T0 = 32'h738631a;
    61: T0 = 32'h60789f2d;
    62: T0 = 32'h4c23519e;
    63: T0 = 32'hf63c6b8b;
    64: T0 = 32'h1be4b25d;
    65: T0 = 32'h4b22709d;
    66: T0 = 32'h68be5f3c;
    67: T0 = 32'h96fc32e;
    68: T0 = 32'h1334340a;
    69: T0 = 32'ha68b9887;
    70: T0 = 32'hd52ff779;
    71: T0 = 32'ha3718539;
    72: T0 = 32'h8e32ad8f;
    73: T0 = 32'he087a07e;
    74: T0 = 32'h7934a723;
    75: T0 = 32'h4d51f90b;
    76: T0 = 32'h556e89af;
    77: T0 = 32'h6a6cf6ce;
    78: T0 = 32'h949ac2c1;
    79: T0 = 32'h539a49f4;
    80: T0 = 32'h67a26f5b;
    81: T0 = 32'h199b0f74;
    82: T0 = 32'h771923ed;
    83: T0 = 32'hbd1ec795;
    84: T0 = 32'h3aba6e5;
    85: T0 = 32'he783a523;
    86: T0 = 32'hdfaf3d00;
    87: T0 = 32'h6ed53e6f;
    88: T0 = 32'ha89a1904;
    89: T0 = 32'h7fc91f49;
    90: T0 = 32'ha3d27fb1;
    91: T0 = 32'he54d7946;
    92: T0 = 32'hb627bec6;
    93: T0 = 32'hb218b3cd;
    94: T0 = 32'hdf430d37;
    95: T0 = 32'hd89c668f;
    96: T0 = 32'h48cbe995;
    97: T0 = 32'he2469760;
    98: T0 = 32'hb2fc4093;
    99: T0 = 32'he6c09ed5;
    100: T0 = 32'h7ef7ddf5;
    101: T0 = 32'h6e350f70;
    102: T0 = 32'h67cce46;
    103: T0 = 32'h5822e9dd;
    104: T0 = 32'h77255769;
    105: T0 = 32'h8c366883;
    106: T0 = 32'h5f29a2d9;
    107: T0 = 32'h5bf022f0;
    108: T0 = 32'h59d65b49;
    109: T0 = 32'h57e73b75;
    110: T0 = 32'h261539f8;
    111: T0 = 32'hb9cf3e5b;
    112: T0 = 32'h23166883;
    113: T0 = 32'h8599975a;
    114: T0 = 32'h1ec3340e;
    115: T0 = 32'h54bf1eef;
    116: T0 = 32'hfa55b573;
    117: T0 = 32'h99eb1e37;
    118: T0 = 32'h5b234681;
    119: T0 = 32'hce213f93;
    120: T0 = 32'hf0c41b19;
    121: T0 = 32'h5c6b00ca;
    122: T0 = 32'h449436e0;
    123: T0 = 32'h907bc3b5;
    124: T0 = 32'h3a71bf81;
    125: T0 = 32'h114afb43;
    126: T0 = 32'h69738981;
    127: T0 = 32'h7b650c19;
    128: T0 = 32'hbc45b3a1;
    129: T0 = 32'hfe431cab;
    130: T0 = 32'h90e96812;
    131: T0 = 32'h58fcb6ec;
    132: T0 = 32'h456c0ade;
    133: T0 = 32'h3e001894;
    134: T0 = 32'h8826bee6;
    135: T0 = 32'h5519e095;
    136: T0 = 32'hb7296753;
    137: T0 = 32'ha59cb501;
    138: T0 = 32'h5a2944b9;
    139: T0 = 32'h3aa39bca;
    140: T0 = 32'h98e70990;
    141: T0 = 32'h89af0977;
    142: T0 = 32'h3389f48f;
    143: T0 = 32'hb43f945;
    144: T0 = 32'h35986b04;
    145: T0 = 32'h7a170a2c;
    146: T0 = 32'h355869f9;
    147: T0 = 32'h79f40114;
    148: T0 = 32'h97263fc5;
    149: T0 = 32'h2784b42c;
    150: T0 = 32'hbb06b344;
    151: T0 = 32'h3fd60d7f;
    152: T0 = 32'hd7e97d0d;
    153: T0 = 32'h7f0c7840;
    154: T0 = 32'h22d10285;
    155: T0 = 32'he3a92be6;
    156: T0 = 32'hbac4a809;
    157: T0 = 32'h9b833eac;
    158: T0 = 32'hbad51d9b;
    159: T0 = 32'h2dd92738;
    160: T0 = 32'h2c59e753;
    161: T0 = 32'h63468b76;
    162: T0 = 32'hf2ec2377;
    163: T0 = 32'h8643efd3;
    164: T0 = 32'h6cf53f25;
    165: T0 = 32'h6eb9e441;
    166: T0 = 32'h263cbd00;
    167: T0 = 32'h505ffe4d;
    168: T0 = 32'h37221d25;
    169: T0 = 32'h98945e49;
    170: T0 = 32'h7d0f3bb5;
    171: T0 = 32'h57d47156;
    172: T0 = 32'h54dcb2d6;
    173: T0 = 32'h7777b38c;
    174: T0 = 32'h64b44d37;
    175: T0 = 32'h318b2682;
    176: T0 = 32'ha736d08b;
    177: T0 = 32'h5a5e37fa;
    178: T0 = 32'haf1c274c;
    179: T0 = 32'haf684693;
    180: T0 = 32'h5b2ea85;
    181: T0 = 32'h66040fe5;
    182: T0 = 32'ha4c46cb4;
    183: T0 = 32'hb1d83b0c;
    184: T0 = 32'h1e2acc20;
    185: T0 = 32'h398c399c;
    186: T0 = 32'hbb5b9608;
    187: T0 = 32'hef8462d1;
    188: T0 = 32'h41c67f6b;
    189: T0 = 32'he6f6268d;
    190: T0 = 32'h96a8718d;
    191: T0 = 32'he49c4a56;
    192: T0 = 32'he7aa49d9;
    193: T0 = 32'h6f6ac622;
    194: T0 = 32'h6844860b;
    195: T0 = 32'h9bae21b;
    196: T0 = 32'h5175eeb5;
    197: T0 = 32'hbe437758;
    198: T0 = 32'h9926ec0e;
    199: T0 = 32'hba11088e;
    200: T0 = 32'h9e795b88;
    201: T0 = 32'h65553fa3;
    202: T0 = 32'hf451ed44;
    203: T0 = 32'h39d12731;
    204: T0 = 32'hb76f250;
    205: T0 = 32'he8486d64;
    206: T0 = 32'h97dada2e;
    207: T0 = 32'h21d90fba;
    208: T0 = 32'h272b4d58;
    209: T0 = 32'h9ce350cf;
    210: T0 = 32'hb8f38d9e;
    211: T0 = 32'h76f5417f;
    212: T0 = 32'hfee9de0a;
    213: T0 = 32'hb970f93f;
    214: T0 = 32'hc342e439;
    215: T0 = 32'h5dabbc88;
    216: T0 = 32'h77c0cccd;
    217: T0 = 32'hb032e8f6;
    218: T0 = 32'hce898b47;
    219: T0 = 32'h3b3b3c3f;
    220: T0 = 32'hf885013f;
    221: T0 = 32'h95efe6ca;
    222: T0 = 32'h538f5383;
    223: T0 = 32'h2b6305b0;
    224: T0 = 32'h104ca610;
    225: T0 = 32'hef7550e7;
    226: T0 = 32'h4a5c817a;
    227: T0 = 32'h9ff227d;
    228: T0 = 32'h8154da7b;
    229: T0 = 32'h3347593d;
    230: T0 = 32'hb883e375;
    231: T0 = 32'hbf40ab1a;
    232: T0 = 32'hdc6f80c7;
    233: T0 = 32'h75476836;
    234: T0 = 32'h78740440;
    235: T0 = 32'hba90553f;
    236: T0 = 32'h7b766dbc;
    237: T0 = 32'h8c06c33;
    238: T0 = 32'hbf9892b6;
    239: T0 = 32'h7d9913b4;
    240: T0 = 32'h77a850d9;
    241: T0 = 32'h108d578f;
    242: T0 = 32'hf59b17ae;
    243: T0 = 32'hff8346eb;
    244: T0 = 32'h9e8adfc8;
    245: T0 = 32'h619d47b5;
    246: T0 = 32'hfedae4dd;
    247: T0 = 32'ha0e62b18;
    248: T0 = 32'hc1b4db88;
    249: T0 = 32'hfa7b23fe;
    250: T0 = 32'ha704964f;
    251: T0 = 32'hc13cf41b;
    252: T0 = 32'h9689133c;
    253: T0 = 32'h56b5ed49;
    254: T0 = 32'h44741364;
    255: T0 = 32'hf6cecd93;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[7:0];
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T6 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_21(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[7:0] T5;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T6;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (T5)
    0: T0 = 32'hebe4f012;
    1: T0 = 32'h17eca35a;
    2: T0 = 32'hebb3ae4e;
    3: T0 = 32'ha28106e6;
    4: T0 = 32'hfc12e626;
    5: T0 = 32'h430c4e26;
    6: T0 = 32'he6c039ca;
    7: T0 = 32'hbcaeab1e;
    8: T0 = 32'h1a643b07;
    9: T0 = 32'h13fa13cb;
    10: T0 = 32'hbfc9efe1;
    11: T0 = 32'h7d37d107;
    12: T0 = 32'h45c2f825;
    13: T0 = 32'hf25ef2c9;
    14: T0 = 32'h16ac0d11;
    15: T0 = 32'hee3e0cde;
    16: T0 = 32'he3e710aa;
    17: T0 = 32'ha720f5ab;
    18: T0 = 32'h88e5f642;
    19: T0 = 32'hc07376ab;
    20: T0 = 32'h255c8f8;
    21: T0 = 32'hbafbcfbc;
    22: T0 = 32'h112d499f;
    23: T0 = 32'he0446390;
    24: T0 = 32'h2c5383fa;
    25: T0 = 32'h845818b;
    26: T0 = 32'h7c26514c;
    27: T0 = 32'h1cc5c419;
    28: T0 = 32'h17f43337;
    29: T0 = 32'h5c884045;
    30: T0 = 32'h2cbb6bce;
    31: T0 = 32'h11fa8957;
    32: T0 = 32'hf7047852;
    33: T0 = 32'h90dbe43c;
    34: T0 = 32'h5793964a;
    35: T0 = 32'h578e20ba;
    36: T0 = 32'h2ebe6f1;
    37: T0 = 32'hdfc8169d;
    38: T0 = 32'hc5b5e05f;
    39: T0 = 32'h64dd0f9a;
    40: T0 = 32'h31184b9c;
    41: T0 = 32'hdb883bea;
    42: T0 = 32'h22fe67c4;
    43: T0 = 32'h866727b7;
    44: T0 = 32'hb419e6b5;
    45: T0 = 32'h333f7626;
    46: T0 = 32'hef499eba;
    47: T0 = 32'hd3641f3a;
    48: T0 = 32'hccc34943;
    49: T0 = 32'ha2058760;
    50: T0 = 32'h13fd2643;
    51: T0 = 32'h4d3e2cd0;
    52: T0 = 32'hb4effb4;
    53: T0 = 32'h3eeae744;
    54: T0 = 32'h181d1c44;
    55: T0 = 32'hf6513d8f;
    56: T0 = 32'he51b5f2c;
    57: T0 = 32'h2d953a8b;
    58: T0 = 32'h90267e85;
    59: T0 = 32'h4ea65a4;
    60: T0 = 32'hb39fb3cf;
    61: T0 = 32'hda13aac;
    62: T0 = 32'heb530d2e;
    63: T0 = 32'h90c5269b;
    64: T0 = 32'h18945dcf;
    65: T0 = 32'ha4aae832;
    66: T0 = 32'h78e7c2c1;
    67: T0 = 32'h80126832;
    68: T0 = 32'he27d429c;
    69: T0 = 32'hda7be7c0;
    70: T0 = 32'h492d34be;
    71: T0 = 32'h46b51aac;
    72: T0 = 32'he2d4d9f8;
    73: T0 = 32'hc153bf2b;
    74: T0 = 32'hfc2e7f3f;
    75: T0 = 32'h14f64c2;
    76: T0 = 32'h5e5a727e;
    77: T0 = 32'h41381625;
    78: T0 = 32'hc33ee2e;
    79: T0 = 32'h535a63aa;
    80: T0 = 32'hfb66a4b1;
    81: T0 = 32'h10bd1ecb;
    82: T0 = 32'hd5b9703c;
    83: T0 = 32'h5d3bbeed;
    84: T0 = 32'h380a9bfb;
    85: T0 = 32'h418e1927;
    86: T0 = 32'h7adb4bc1;
    87: T0 = 32'he17ff0dd;
    88: T0 = 32'h89b62663;
    89: T0 = 32'h22db5085;
    90: T0 = 32'h85f6064b;
    91: T0 = 32'hc57a1a19;
    92: T0 = 32'hbe8b0d28;
    93: T0 = 32'h54a56d73;
    94: T0 = 32'h4d46316d;
    95: T0 = 32'hd6a09c47;
    96: T0 = 32'hd9f55b87;
    97: T0 = 32'hee11155c;
    98: T0 = 32'h8a6479f4;
    99: T0 = 32'h40239784;
    100: T0 = 32'hb65727c4;
    101: T0 = 32'hf4f7b686;
    102: T0 = 32'h15355bc0;
    103: T0 = 32'hc244e77d;
    104: T0 = 32'h6cd73f28;
    105: T0 = 32'h594900d0;
    106: T0 = 32'h7c02a0ab;
    107: T0 = 32'h6c8bae2;
    108: T0 = 32'h27f49b03;
    109: T0 = 32'hecc0badc;
    110: T0 = 32'h2f3529c9;
    111: T0 = 32'h553ea45b;
    112: T0 = 32'h3e00fa5f;
    113: T0 = 32'h70a47198;
    114: T0 = 32'h352a1fbc;
    115: T0 = 32'h3403492a;
    116: T0 = 32'hbe8c0308;
    117: T0 = 32'he3bfaa8f;
    118: T0 = 32'h56def739;
    119: T0 = 32'haee9320;
    120: T0 = 32'h48b7ec92;
    121: T0 = 32'h767281fc;
    122: T0 = 32'ha389ab22;
    123: T0 = 32'h44d8d90b;
    124: T0 = 32'h87d084a7;
    125: T0 = 32'h7e80d1c8;
    126: T0 = 32'h4876a2c1;
    127: T0 = 32'hbc9c11b9;
    128: T0 = 32'hb85fcf49;
    129: T0 = 32'hef5bca35;
    130: T0 = 32'hbf4c451;
    131: T0 = 32'h22ff6a53;
    132: T0 = 32'hed137af5;
    133: T0 = 32'hbe75a5c0;
    134: T0 = 32'he421f404;
    135: T0 = 32'h9c083e4d;
    136: T0 = 32'hfe4fc9ec;
    137: T0 = 32'h5d2ffe2a;
    138: T0 = 32'h1e491ec5;
    139: T0 = 32'hbb932cf7;
    140: T0 = 32'h7944fb5e;
    141: T0 = 32'hba567ea5;
    142: T0 = 32'hbba8842a;
    143: T0 = 32'h4931736a;
    144: T0 = 32'h668a59db;
    145: T0 = 32'h6306d758;
    146: T0 = 32'he2eeae4b;
    147: T0 = 32'h874346da;
    148: T0 = 32'h24f5ee85;
    149: T0 = 32'hceb947b1;
    150: T0 = 32'h173c6c94;
    151: T0 = 32'h30552a9f;
    152: T0 = 32'h1a265b08;
    153: T0 = 32'h88853bda;
    154: T0 = 32'h5b27e7cd;
    155: T0 = 32'h9f44e636;
    156: T0 = 32'h51bdf21a;
    157: T0 = 32'h77b73665;
    158: T0 = 32'h64b0ddbe;
    159: T0 = 32'h11a36e1b;
    160: T0 = 32'hb716b664;
    161: T0 = 32'h6346d0b1;
    162: T0 = 32'ha2ec6cb1;
    163: T0 = 32'h86c2b85c;
    164: T0 = 32'h20fd003c;
    165: T0 = 32'hfef102d8;
    166: T0 = 32'h63cda6a;
    167: T0 = 32'h505545b7;
    168: T0 = 32'h172314f2;
    169: T0 = 32'h8884dd27;
    170: T0 = 32'h792e48b2;
    171: T0 = 32'h83c4399b;
    172: T0 = 32'h51df84a5;
    173: T0 = 32'h7ea74936;
    174: T0 = 32'h2eb0a4e3;
    175: T0 = 32'h108b9935;
    176: T0 = 32'h27367e76;
    177: T0 = 32'h8f08cf14;
    178: T0 = 32'h98452241;
    179: T0 = 32'h61f10d8a;
    180: T0 = 32'hf7556517;
    181: T0 = 32'h19dd7ceb;
    182: T0 = 32'hb16bbd62;
    183: T0 = 32'hca041e7f;
    184: T0 = 32'hf6c5563e;
    185: T0 = 32'hec65075d;
    186: T0 = 32'h6e40ee56;
    187: T0 = 32'hb89d4156;
    188: T0 = 32'ha646eb4;
    189: T0 = 32'h5d5abfe8;
    190: T0 = 32'hbcbd9c39;
    191: T0 = 32'h39fc4eab;
    192: T0 = 32'h320c8bbc;
    193: T0 = 32'haf895d89;
    194: T0 = 32'hc4d79bc;
    195: T0 = 32'h49bf99ad;
    196: T0 = 32'h9355814a;
    197: T0 = 32'h996fa8a7;
    198: T0 = 32'h1b376773;
    199: T0 = 32'hea44c1b0;
    200: T0 = 32'he4c566d3;
    201: T0 = 32'hf56d81f4;
    202: T0 = 32'h2c04a83b;
    203: T0 = 32'h90599a09;
    204: T0 = 32'h2e7805a8;
    205: T0 = 32'h5908d8d2;
    206: T0 = 32'h2b37b2d1;
    207: T0 = 32'h79ddd165;
    208: T0 = 32'hae44cf7a;
    209: T0 = 32'h509fe8e7;
    210: T0 = 32'h37da82d2;
    211: T0 = 32'hbb6c78f5;
    212: T0 = 32'h7afdaf3;
    213: T0 = 32'h6f898134;
    214: T0 = 32'h5f278224;
    215: T0 = 32'h629476ce;
    216: T0 = 32'h2b38c4f6;
    217: T0 = 32'hef00fe24;
    218: T0 = 32'h339a1a5f;
    219: T0 = 32'ha7ed0576;
    220: T0 = 32'hf287607a;
    221: T0 = 32'hbf330d38;
    222: T0 = 32'ha7497332;
    223: T0 = 32'h518db326;
    224: T0 = 32'h4d978532;
    225: T0 = 32'h2264faeb;
    226: T0 = 32'hb06954be;
    227: T0 = 32'h7400fae5;
    228: T0 = 32'hf8acdafa;
    229: T0 = 32'h407ac93f;
    230: T0 = 32'h8a1e72f9;
    231: T0 = 32'h5b797290;
    232: T0 = 32'h579180c3;
    233: T0 = 32'ha0d2c5b4;
    234: T0 = 32'hc881095f;
    235: T0 = 32'h41ba181b;
    236: T0 = 32'h9b89113e;
    237: T0 = 32'h85854471;
    238: T0 = 32'h5a126343;
    239: T0 = 32'ha8c3f1c6;
    240: T0 = 32'h9175346c;
    241: T0 = 32'h967ae8b4;
    242: T0 = 32'h68e58e00;
    243: T0 = 32'hcaf118ba;
    244: T0 = 32'ha930420f;
    245: T0 = 32'h581d8dbd;
    246: T0 = 32'ha8ed36f6;
    247: T0 = 32'h3430c412;
    248: T0 = 32'h94e8a5f8;
    249: T0 = 32'hc4f6ff6e;
    250: T0 = 32'hff74458f;
    251: T0 = 32'hdb1655ca;
    252: T0 = 32'h784e6238;
    253: T0 = 32'h207e0512;
    254: T0 = 32'h8caad6dc;
    255: T0 = 32'h5675eb26;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[7:0];
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T6 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_22(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[7:0] T5;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T6;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (T5)
    0: T0 = 32'h3fba80b8;
    1: T0 = 32'h9abd25cb;
    2: T0 = 32'h1d10fefd;
    3: T0 = 32'h78b596a6;
    4: T0 = 32'hd92a9d4a;
    5: T0 = 32'h9142cb63;
    6: T0 = 32'hc9c331e2;
    7: T0 = 32'hefa0b328;
    8: T0 = 32'hc5d9ba27;
    9: T0 = 32'h777a80fd;
    10: T0 = 32'ha6d0fb63;
    11: T0 = 32'h7833d85e;
    12: T0 = 32'hbe069d69;
    13: T0 = 32'h81c8f6db;
    14: T0 = 32'h9b4f0751;
    15: T0 = 32'hec7485d5;
    16: T0 = 32'h58c9fcdd;
    17: T0 = 32'h85da8f76;
    18: T0 = 32'hc7432241;
    19: T0 = 32'h33cbecd3;
    20: T0 = 32'h614165b5;
    21: T0 = 32'hfd724651;
    22: T0 = 32'h63700d0a;
    23: T0 = 32'h8dac7e0f;
    24: T0 = 32'h1b4e1f3c;
    25: T0 = 32'h9a37078b;
    26: T0 = 32'had93e92;
    27: T0 = 32'hba706954;
    28: T0 = 32'h4534b6c6;
    29: T0 = 32'hf5c73be5;
    30: T0 = 32'hf2e90d2c;
    31: T0 = 32'hb264ecb;
    32: T0 = 32'h16df6b24;
    33: T0 = 32'h408f902c;
    34: T0 = 32'h35ca4970;
    35: T0 = 32'he2d57154;
    36: T0 = 32'hd7f13950;
    37: T0 = 32'h699db29e;
    38: T0 = 32'hf43d21b;
    39: T0 = 32'hc265de9;
    40: T0 = 32'h7344e0dc;
    41: T0 = 32'hfe2afca4;
    42: T0 = 32'ha80930b9;
    43: T0 = 32'hf0d82be4;
    44: T0 = 32'h6ed148c3;
    45: T0 = 32'h7b7f38ae;
    46: T0 = 32'h1a1fa09b;
    47: T0 = 32'ha9cc3338;
    48: T0 = 32'hea5c9eb9;
    49: T0 = 32'h9dd94d13;
    50: T0 = 32'h5b1779b5;
    51: T0 = 32'h8f1b9b0a;
    52: T0 = 32'h5a0b1146;
    53: T0 = 32'hc285f8c3;
    54: T0 = 32'hf5f18f8a;
    55: T0 = 32'ha406c0d5;
    56: T0 = 32'ha8b6777a;
    57: T0 = 32'h49e886d0;
    58: T0 = 32'ha3f22c33;
    59: T0 = 32'h855fab68;
    60: T0 = 32'h66798888;
    61: T0 = 32'h721edd5b;
    62: T0 = 32'hcd65ce70;
    63: T0 = 32'hd634d8c9;
    64: T0 = 32'h79cb7b22;
    65: T0 = 32'hac30f0b8;
    66: T0 = 32'h7c511c6c;
    67: T0 = 32'h51b494ac;
    68: T0 = 32'hbae4a60a;
    69: T0 = 32'h947a0c3f;
    70: T0 = 32'h991f33f9;
    71: T0 = 32'hc3d1cf33;
    72: T0 = 32'he4d32082;
    73: T0 = 32'h235bd1ed;
    74: T0 = 32'hc4d06683;
    75: T0 = 32'hac7b894e;
    76: T0 = 32'h9b68abac;
    77: T0 = 32'hc9881516;
    78: T0 = 32'h99db8793;
    79: T0 = 32'hbf4ed9a;
    80: T0 = 32'hf86d83bd;
    81: T0 = 32'h8198c503;
    82: T0 = 32'hd8b71b7;
    83: T0 = 32'hf18fb045;
    84: T0 = 32'h8780196a;
    85: T0 = 32'h9acc30c2;
    86: T0 = 32'hf7738626;
    87: T0 = 32'h32e550e5;
    88: T0 = 32'h28a0f2fb;
    89: T0 = 32'hfecbecb4;
    90: T0 = 32'ha1d418d9;
    91: T0 = 32'h980d86f0;
    92: T0 = 32'h846a6849;
    93: T0 = 32'h737808be;
    94: T0 = 32'h8cf8f2ba;
    95: T0 = 32'h43dab378;
    96: T0 = 32'he0d3ec53;
    97: T0 = 32'haf601274;
    98: T0 = 32'hc8236064;
    99: T0 = 32'hc4932eef;
    100: T0 = 32'hb850ffc1;
    101: T0 = 32'h47a0135;
    102: T0 = 32'ha0584ac5;
    103: T0 = 32'h8d6b2d9f;
    104: T0 = 32'hd4c67f0c;
    105: T0 = 32'h10f63002;
    106: T0 = 32'hce65a6a4;
    107: T0 = 32'h5896bb95;
    108: T0 = 32'h5e89d81;
    109: T0 = 32'he4d4bb41;
    110: T0 = 32'h18b6192a;
    111: T0 = 32'haeb20e1f;
    112: T0 = 32'hb2e8f7dd;
    113: T0 = 32'h94c3cb16;
    114: T0 = 32'ha6e3ef93;
    115: T0 = 32'h9642f912;
    116: T0 = 32'heed1210c;
    117: T0 = 32'hccbcf4c0;
    118: T0 = 32'hc774b42a;
    119: T0 = 32'hc8fd8a7;
    120: T0 = 32'h7a4c39b8;
    121: T0 = 32'h9b229f6e;
    122: T0 = 32'hf8bf932;
    123: T0 = 32'h4f5f7552;
    124: T0 = 32'hdc9156de;
    125: T0 = 32'hb37ed58c;
    126: T0 = 32'h5265f634;
    127: T0 = 32'h4b665be9;
    128: T0 = 32'haccfb67e;
    129: T0 = 32'h794768d5;
    130: T0 = 32'h8f3c6375;
    131: T0 = 32'h3e638975;
    132: T0 = 32'h8e863a0b;
    133: T0 = 32'h269458af;
    134: T0 = 32'ha410b1f8;
    135: T0 = 32'h6bc4b675;
    136: T0 = 32'h6d6f24d7;
    137: T0 = 32'h1b08d174;
    138: T0 = 32'h170b8b32;
    139: T0 = 32'h77a8595e;
    140: T0 = 32'he3c50cb4;
    141: T0 = 32'h9a438c9b;
    142: T0 = 32'h3b555675;
    143: T0 = 32'h92bc3c4;
    144: T0 = 32'h240ba664;
    145: T0 = 32'h7b4d8141;
    146: T0 = 32'he11475b4;
    147: T0 = 32'h2fc9b9c5;
    148: T0 = 32'h2112157a;
    149: T0 = 32'h67046ada;
    150: T0 = 32'ha6c81b6b;
    151: T0 = 32'hf51ed3e5;
    152: T0 = 32'h1d263237;
    153: T0 = 32'hc9bc4e85;
    154: T0 = 32'hbf6a58b2;
    155: T0 = 32'h7b269989;
    156: T0 = 32'h65e78cc5;
    157: T0 = 32'hf2d778fa;
    158: T0 = 32'h90acae63;
    159: T0 = 32'he4b39434;
    160: T0 = 32'h73b85dee;
    161: T0 = 32'h97cded33;
    162: T0 = 32'h4983b643;
    163: T0 = 32'h7bfd7d92;
    164: T0 = 32'hc310410c;
    165: T0 = 32'h1b8ce4d2;
    166: T0 = 32'hacc2383e;
    167: T0 = 32'h9c2e5a26;
    168: T0 = 32'hf4e592ba;
    169: T0 = 32'hfcbea7ed;
    170: T0 = 32'hb9757915;
    171: T0 = 32'h383bc4c2;
    172: T0 = 32'h28e6727e;
    173: T0 = 32'h934fd0ac;
    174: T0 = 32'h949cee2e;
    175: T0 = 32'h6853f1e9;
    176: T0 = 32'h61603094;
    177: T0 = 32'h50953719;
    178: T0 = 32'h15983f06;
    179: T0 = 32'h6d1f95ce;
    180: T0 = 32'h930e6182;
    181: T0 = 32'h618d1a8f;
    182: T0 = 32'h5edb09ca;
    183: T0 = 32'hd07eab95;
    184: T0 = 32'h81353773;
    185: T0 = 32'h7c09019b;
    186: T0 = 32'ha176e1a8;
    187: T0 = 32'hc4289811;
    188: T0 = 32'h3fab8e85;
    189: T0 = 32'h1e91c056;
    190: T0 = 32'he907bc8d;
    191: T0 = 32'hf48c9857;
    192: T0 = 32'hcad56f75;
    193: T0 = 32'h32b64ad4;
    194: T0 = 32'h375909fd;
    195: T0 = 32'h7fac8156;
    196: T0 = 32'h9faf3467;
    197: T0 = 32'h21093ca3;
    198: T0 = 32'h5aafa560;
    199: T0 = 32'h4beb8c3f;
    200: T0 = 32'he334642f;
    201: T0 = 32'h37737254;
    202: T0 = 32'h1d19ef3;
    203: T0 = 32'he1a8016e;
    204: T0 = 32'hdb012eac;
    205: T0 = 32'h8c91ab88;
    206: T0 = 32'hc152f711;
    207: T0 = 32'hbe8566a0;
    208: T0 = 32'h4c5d6b2c;
    209: T0 = 32'hbe26708c;
    210: T0 = 32'ha864810a;
    211: T0 = 32'h68d10174;
    212: T0 = 32'h3914f04a;
    213: T0 = 32'h2636be9c;
    214: T0 = 32'h30d8e275;
    215: T0 = 32'h1b621db2;
    216: T0 = 32'hc6ffe0d1;
    217: T0 = 32'h7777f874;
    218: T0 = 32'hbd0554c8;
    219: T0 = 32'h78bb87ab;
    220: T0 = 32'h4be66aa9;
    221: T0 = 32'hedc18cbe;
    222: T0 = 32'h12bef69a;
    223: T0 = 32'hbcd31330;
    224: T0 = 32'h726d0928;
    225: T0 = 32'h1aebe8ab;
    226: T0 = 32'h2d70864a;
    227: T0 = 32'h397d6070;
    228: T0 = 32'hd72adafb;
    229: T0 = 32'h2500c5dc;
    230: T0 = 32'hb80ae03d;
    231: T0 = 32'hbd90180a;
    232: T0 = 32'h8cd980d2;
    233: T0 = 32'h7714fda6;
    234: T0 = 32'h25d95c5d;
    235: T0 = 32'heaab443f;
    236: T0 = 32'hff46637d;
    237: T0 = 32'h88094c24;
    238: T0 = 32'h9b4fc2a2;
    239: T0 = 32'hddc33a2;
    240: T0 = 32'h4c49ef0a;
    241: T0 = 32'h4de10e6c;
    242: T0 = 32'hf2a3216a;
    243: T0 = 32'h9403e7b5;
    244: T0 = 32'h38dbbef1;
    245: T0 = 32'hecf0a524;
    246: T0 = 32'h67943c80;
    247: T0 = 32'hc41fbe4b;
    248: T0 = 32'h288edf24;
    249: T0 = 32'h93c87e59;
    250: T0 = 32'hfaf7bc1;
    251: T0 = 32'h555cc1f6;
    252: T0 = 32'h5b1bb4e;
    253: T0 = 32'h6259b2f8;
    254: T0 = 32'h4e24399b;
    255: T0 = 32'hd626278b;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[7:0];
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T6 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_23(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[7:0] T5;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T6;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (T5)
    0: T0 = 32'hc9655dfa;
    1: T0 = 32'h19d9ec43;
    2: T0 = 32'h7d39b2c1;
    3: T0 = 32'h8d1a6e93;
    4: T0 = 32'h42abcd14;
    5: T0 = 32'hdbcae761;
    6: T0 = 32'hd9a50dae;
    7: T0 = 32'he7953ace;
    8: T0 = 32'h807293ae;
    9: T0 = 32'hcbc90afb;
    10: T0 = 32'ha2f2fb57;
    11: T0 = 32'ha44d4425;
    12: T0 = 32'hb631f37f;
    13: T0 = 32'h7318f4a1;
    14: T0 = 32'hed424f24;
    15: T0 = 32'h589c27cb;
    16: T0 = 32'he92f87aa;
    17: T0 = 32'h50720949;
    18: T0 = 32'h629a79fd;
    19: T0 = 32'h974cc711;
    20: T0 = 32'h93a19cc;
    21: T0 = 32'he608a962;
    22: T0 = 32'h6d9d1e20;
    23: T0 = 32'h75f9f6e9;
    24: T0 = 32'h8b3aec67;
    25: T0 = 32'h192e858;
    26: T0 = 32'h8b7c18af;
    27: T0 = 32'he576a8ec;
    28: T0 = 32'hd10b994a;
    29: T0 = 32'h223da899;
    30: T0 = 32'hc50829db;
    31: T0 = 32'hc603e045;
    32: T0 = 32'h5dbe91db;
    33: T0 = 32'h6a63f58b;
    34: T0 = 32'h9074964a;
    35: T0 = 32'h7c64c6ab;
    36: T0 = 32'h7ceccad9;
    37: T0 = 32'h7cf2c765;
    38: T0 = 32'h21c69b5;
    39: T0 = 32'h5919a284;
    40: T0 = 32'h671b8b88;
    41: T0 = 32'hb516a79d;
    42: T0 = 32'h4c89dd4d;
    43: T0 = 32'h26a8c41b;
    44: T0 = 32'he885737e;
    45: T0 = 32'h8d874471;
    46: T0 = 32'h7b01530e;
    47: T0 = 32'h29ebc8cf;
    48: T0 = 32'h1e1a845d;
    49: T0 = 32'h976e0755;
    50: T0 = 32'h2dd97ffd;
    51: T0 = 32'hebfdcfc6;
    52: T0 = 32'hdf003d0d;
    53: T0 = 32'h2b0c6843;
    54: T0 = 32'hb5e35d02;
    55: T0 = 32'h3d22b06d;
    56: T0 = 32'hb66d5f25;
    57: T0 = 32'hf62e065a;
    58: T0 = 32'hb759baa2;
    59: T0 = 32'hf9b77b15;
    60: T0 = 32'hd8469cc3;
    61: T0 = 32'hbb5ebbcd;
    62: T0 = 32'h84dc5965;
    63: T0 = 32'h6d598c55;
    64: T0 = 32'he1c5a2b0;
    65: T0 = 32'hc4f025c9;
    66: T0 = 32'hffc379bc;
    67: T0 = 32'h168b85ed;
    68: T0 = 32'hfeeb184a;
    69: T0 = 32'hd83a9aaf;
    70: T0 = 32'h4ff331fb;
    71: T0 = 32'h4dbbb328;
    72: T0 = 32'hfb00b687;
    73: T0 = 32'h92ea80f5;
    74: T0 = 32'h85bd8ba3;
    75: T0 = 32'hdf5fd81f;
    76: T0 = 32'ha0199d25;
    77: T0 = 32'h637cc0db;
    78: T0 = 32'hc0211bd1;
    79: T0 = 32'he62781d5;
    80: T0 = 32'hd9d5957f;
    81: T0 = 32'h118e68e5;
    82: T0 = 32'hb429cad1;
    83: T0 = 32'hff00e991;
    84: T0 = 32'h7eadc83d;
    85: T0 = 32'h8b99804d;
    86: T0 = 32'h939c3436;
    87: T0 = 32'h5297f26c;
    88: T0 = 32'h7761c4f2;
    89: T0 = 32'he350ff6c;
    90: T0 = 32'hb7b85b1f;
    91: T0 = 32'h518c184a;
    92: T0 = 32'hda83217e;
    93: T0 = 32'h511b0c8b;
    94: T0 = 32'h44547275;
    95: T0 = 32'hf0cffbe4;
    96: T0 = 32'h993f828f;
    97: T0 = 32'h6805256a;
    98: T0 = 32'hd0366ac5;
    99: T0 = 32'h402ded1;
    100: T0 = 32'h287e618d;
    101: T0 = 32'hf6724f43;
    102: T0 = 32'h529c0c06;
    103: T0 = 32'hc25f7245;
    104: T0 = 32'h2912fe2e;
    105: T0 = 32'h991ac0d;
    106: T0 = 32'h4fa6f37d;
    107: T0 = 32'h86406ed0;
    108: T0 = 32'h25b91f5b;
    109: T0 = 32'h66a51a35;
    110: T0 = 32'h69252ddc;
    111: T0 = 32'h86a6ca5d;
    112: T0 = 32'h1f3a5f5b;
    113: T0 = 32'h78927f1c;
    114: T0 = 32'h67da893e;
    115: T0 = 32'hbf4e4133;
    116: T0 = 32'h6aab6c2;
    117: T0 = 32'hce8bbda7;
    118: T0 = 32'h4f2fe655;
    119: T0 = 32'h21f18c7a;
    120: T0 = 32'h8b9a6fcd;
    121: T0 = 32'hf0ee2f2;
    122: T0 = 32'h33daa6c3;
    123: T0 = 32'he7453776;
    124: T0 = 32'hd11f2208;
    125: T0 = 32'hba3cbfc8;
    126: T0 = 32'hf74340bc;
    127: T0 = 32'hd70c63aa;
    128: T0 = 32'hcd9f8338;
    129: T0 = 32'h68857009;
    130: T0 = 32'h171c593a;
    131: T0 = 32'h3d169174;
    132: T0 = 32'h1fee9afa;
    133: T0 = 32'h6383b9ac;
    134: T0 = 32'h1e9ee351;
    135: T0 = 32'hcacfc771;
    136: T0 = 32'h6db761d1;
    137: T0 = 32'h7771e8b2;
    138: T0 = 32'h85038049;
    139: T0 = 32'hc6b8b6e3;
    140: T0 = 32'ha3814109;
    141: T0 = 32'h4c85cc72;
    142: T0 = 32'h6957f0da;
    143: T0 = 32'hbc9db93d;
    144: T0 = 32'h58591089;
    145: T0 = 32'he9c9f5bb;
    146: T0 = 32'h1747d606;
    147: T0 = 32'he79020ea;
    148: T0 = 32'h6758d8aa;
    149: T0 = 32'hd9f44b1c;
    150: T0 = 32'h471452fb;
    151: T0 = 32'hce06019a;
    152: T0 = 32'h35ed8888;
    153: T0 = 32'hdf2cc3be;
    154: T0 = 32'h2ed3226e;
    155: T0 = 32'hbaacb419;
    156: T0 = 32'h2eb59725;
    157: T0 = 32'hd5436247;
    158: T0 = 32'h7aad82e6;
    159: T0 = 32'h96e98d4;
    160: T0 = 32'h3619192b;
    161: T0 = 32'ha3b07829;
    162: T0 = 32'h54bc802;
    163: T0 = 32'h793b7131;
    164: T0 = 32'h97c5dab8;
    165: T0 = 32'h197bb59c;
    166: T0 = 32'h192fd63d;
    167: T0 = 32'h8b434472;
    168: T0 = 32'ha353c1d8;
    169: T0 = 32'h3207a9e2;
    170: T0 = 32'h4015450d;
    171: T0 = 32'h8448a6e0;
    172: T0 = 32'h9b3d431a;
    173: T0 = 32'hdd810024;
    174: T0 = 32'he8dbe3de;
    175: T0 = 32'h89d9b368;
    176: T0 = 32'h945501ba;
    177: T0 = 32'ha4926c8b;
    178: T0 = 32'hcf72d9cb;
    179: T0 = 32'h960a0351;
    180: T0 = 32'hbecf98ae;
    181: T0 = 32'hcedff773;
    182: T0 = 32'h453d22e5;
    183: T0 = 32'h28c692e0;
    184: T0 = 32'headfe2cb;
    185: T0 = 32'h1b69a1f4;
    186: T0 = 32'h15cbd94f;
    187: T0 = 32'hcf45447a;
    188: T0 = 32'h571a7378;
    189: T0 = 32'h7b1c84f8;
    190: T0 = 32'he57153da;
    191: T0 = 32'h532ce1c5;
    192: T0 = 32'hcc470520;
    193: T0 = 32'hb76c8a65;
    194: T0 = 32'h8a14c053;
    195: T0 = 32'he9f936d5;
    196: T0 = 32'hd715f5ff;
    197: T0 = 32'h3f075778;
    198: T0 = 32'hb06988c6;
    199: T0 = 32'hbe0420d1;
    200: T0 = 32'hf667c34d;
    201: T0 = 32'h7d25fc83;
    202: T0 = 32'h7f585ed5;
    203: T0 = 32'hf89106fc;
    204: T0 = 32'h63e6f938;
    205: T0 = 32'hd8ca2e37;
    206: T0 = 32'hb7bc1d3e;
    207: T0 = 32'h7d39ee44;
    208: T0 = 32'he60cfe55;
    209: T0 = 32'hc909da16;
    210: T0 = 32'h92670633;
    211: T0 = 32'h909be85f;
    212: T0 = 32'h20502795;
    213: T0 = 32'hddf47499;
    214: T0 = 32'h27548408;
    215: T0 = 32'hd624bcd7;
    216: T0 = 32'h298819b1;
    217: T0 = 32'hdc8c5662;
    218: T0 = 32'he8a69f52;
    219: T0 = 32'h12df7755;
    220: T0 = 32'h26fc6480;
    221: T0 = 32'hf34b2b65;
    222: T0 = 32'h3a34d034;
    223: T0 = 32'hc9fa5f29;
    224: T0 = 32'h3730b6b4;
    225: T0 = 32'h38b0f991;
    226: T0 = 32'hf6ab7694;
    227: T0 = 32'h960ef8af;
    228: T0 = 32'h20eb613a;
    229: T0 = 32'hcce248cb;
    230: T0 = 32'hb1ecb3b;
    231: T0 = 32'h41ffd3d0;
    232: T0 = 32'h2f9820f3;
    233: T0 = 32'ha3cac48d;
    234: T0 = 32'h81aef132;
    235: T0 = 32'h87661b11;
    236: T0 = 32'h9ca90487;
    237: T0 = 32'hd5354153;
    238: T0 = 32'h4242be65;
    239: T0 = 32'h8282d864;
    240: T0 = 32'h197394fc;
    241: T0 = 32'h96fe4f93;
    242: T0 = 32'h759b6281;
    243: T0 = 32'h7fb4fe83;
    244: T0 = 32'hd8af011d;
    245: T0 = 32'h11bc6c0;
    246: T0 = 32'h58eb08a2;
    247: T0 = 32'h4bbbe2c5;
    248: T0 = 32'hd2421272;
    249: T0 = 32'h2273870d;
    250: T0 = 32'hc55cf917;
    251: T0 = 32'he17a4c40;
    252: T0 = 32'hdb115776;
    253: T0 = 32'h4a28575;
    254: T0 = 32'hd1427d6c;
    255: T0 = 32'hf645f847;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[7:0];
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T6 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_24(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[7:0] T5;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T6;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (T5)
    0: T0 = 32'h3e59cd9d;
    1: T0 = 32'haf2d5b87;
    2: T0 = 32'hc835a39b;
    3: T0 = 32'h68b1eb11;
    4: T0 = 32'hf1519bed;
    5: T0 = 32'h197cf5e1;
    6: T0 = 32'ha0d0c424;
    7: T0 = 32'h9e2e70c4;
    8: T0 = 32'h55e7dceb;
    9: T0 = 32'h73a652;
    10: T0 = 32'hce25b85f;
    11: T0 = 32'h38382670;
    12: T0 = 32'h2ae4725a;
    13: T0 = 32'h8cc2a9e9;
    14: T0 = 32'h1abe596e;
    15: T0 = 32'he8e2b2e0;
    16: T0 = 32'h332036ee;
    17: T0 = 32'h80142d32;
    18: T0 = 32'h61c9a343;
    19: T0 = 32'h7dbc2d96;
    20: T0 = 32'h116e61b7;
    21: T0 = 32'h3d0a74c8;
    22: T0 = 32'h9ba7b9c6;
    23: T0 = 32'hb1fb4a5f;
    24: T0 = 32'h93385635;
    25: T0 = 32'hbc87bf1b;
    26: T0 = 32'hf4cb54;
    27: T0 = 32'hbba35f52;
    28: T0 = 32'hd81f6654;
    29: T0 = 32'h9d2507a2;
    30: T0 = 32'hf2dabc3e;
    31: T0 = 32'h251dac7;
    32: T0 = 32'hc5d5e626;
    33: T0 = 32'h22858868;
    34: T0 = 32'h1a9c72e1;
    35: T0 = 32'h693ead54;
    36: T0 = 32'h136e0d36;
    37: T0 = 32'h23cb2048;
    38: T0 = 32'h988f196a;
    39: T0 = 32'hf255de6d;
    40: T0 = 32'hc4b11636;
    41: T0 = 32'h67530e1d;
    42: T0 = 32'hb1007ab2;
    43: T0 = 32'h9849ce;
    44: T0 = 32'hbbfaa4e5;
    45: T0 = 32'hc803aaa;
    46: T0 = 32'h9562df3;
    47: T0 = 32'hb499367c;
    48: T0 = 32'hfa151234;
    49: T0 = 32'hcb80ac08;
    50: T0 = 32'h174ba999;
    51: T0 = 32'h35ff9115;
    52: T0 = 32'hc745010f;
    53: T0 = 32'h3de23ccb;
    54: T0 = 32'hd363b254;
    55: T0 = 32'h49098cf5;
    56: T0 = 32'h3b4d6653;
    57: T0 = 32'h1b07a974;
    58: T0 = 32'h95c89d;
    59: T0 = 32'hb8600fea;
    60: T0 = 32'h8a344ac8;
    61: T0 = 32'hbfc38cb6;
    62: T0 = 32'hfabdf498;
    63: T0 = 32'h2903f379;
    64: T0 = 32'h4795f9c;
    65: T0 = 32'ha65d4f06;
    66: T0 = 32'h5ad5a99b;
    67: T0 = 32'h46b58711;
    68: T0 = 32'h6a5b038d;
    69: T0 = 32'h3e4bbdeb;
    70: T0 = 32'h4807a464;
    71: T0 = 32'hd53988f4;
    72: T0 = 32'hf4497549;
    73: T0 = 32'h8b53174;
    74: T0 = 32'h5c7ecd0d;
    75: T0 = 32'h9b32267a;
    76: T0 = 32'h79556a1a;
    77: T0 = 32'h9cd68dfc;
    78: T0 = 32'h279b759c;
    79: T0 = 32'h161e3cb;
    80: T0 = 32'h53247027;
    81: T0 = 32'h59cceeba;
    82: T0 = 32'h82a41624;
    83: T0 = 32'h2ac10cba;
    84: T0 = 32'h4d10662a;
    85: T0 = 32'h67854a94;
    86: T0 = 32'he6d875d9;
    87: T0 = 32'h5c268f1a;
    88: T0 = 32'h1fa61392;
    89: T0 = 32'hdc2a93ef;
    90: T0 = 32'h7b6e6762;
    91: T0 = 32'hf19df19b;
    92: T0 = 32'h6483a5a5;
    93: T0 = 32'h76774342;
    94: T0 = 32'h36a48603;
    95: T0 = 32'hf48b5daf;
    96: T0 = 32'h66b2c901;
    97: T0 = 32'ha12992a3;
    98: T0 = 32'h5c87548a;
    99: T0 = 32'h4c176170;
    100: T0 = 32'hb045d8f8;
    101: T0 = 32'h985fa73c;
    102: T0 = 32'h91d0c635;
    103: T0 = 32'hce6675e2;
    104: T0 = 32'hc0f5e8cc;
    105: T0 = 32'h667bec84;
    106: T0 = 32'heca434ed;
    107: T0 = 32'h478a6b9;
    108: T0 = 32'hb6f9734b;
    109: T0 = 32'h9807abd;
    110: T0 = 32'h876818a;
    111: T0 = 32'hf0ce3538;
    112: T0 = 32'hbb6488a8;
    113: T0 = 32'h4945f1cb;
    114: T0 = 32'hd11cd498;
    115: T0 = 32'h150bb079;
    116: T0 = 32'h404ad96a;
    117: T0 = 32'h55c04a9e;
    118: T0 = 32'h36dada57;
    119: T0 = 32'hc615e994;
    120: T0 = 32'hda5e7fb;
    121: T0 = 32'h7908a8f6;
    122: T0 = 32'h28f2a00e;
    123: T0 = 32'ha4e88cbb;
    124: T0 = 32'ha6b17939;
    125: T0 = 32'hfac34c33;
    126: T0 = 32'h7b64f2c8;
    127: T0 = 32'h88aa1871;
    128: T0 = 32'h153894ec;
    129: T0 = 32'h7f47cd73;
    130: T0 = 32'hfa34e693;
    131: T0 = 32'h8e10fe83;
    132: T0 = 32'h787b003f;
    133: T0 = 32'h6395eec3;
    134: T0 = 32'hb4d409aa;
    135: T0 = 32'hf615f245;
    136: T0 = 32'h6c373272;
    137: T0 = 32'h69d887cd;
    138: T0 = 32'hfe62f917;
    139: T0 = 32'h5bf5c50;
    140: T0 = 32'h27e255f6;
    141: T0 = 32'h221a5575;
    142: T0 = 32'hb246d64;
    143: T0 = 32'hf03ef8c7;
    144: T0 = 32'h7b2b5178;
    145: T0 = 32'h33b4e8a7;
    146: T0 = 32'h348881cb;
    147: T0 = 32'h59bd2111;
    148: T0 = 32'h972cdaf9;
    149: T0 = 32'h210f65bd;
    150: T0 = 32'hbacba635;
    151: T0 = 32'h73f70ac6;
    152: T0 = 32'h8531c8cb;
    153: T0 = 32'h65c3f926;
    154: T0 = 32'hb1745c5d;
    155: T0 = 32'he1ab247a;
    156: T0 = 32'h9acb7278;
    157: T0 = 32'hab96ca8;
    158: T0 = 32'h8156d21e;
    159: T0 = 32'hb4d92ba2;
    160: T0 = 32'hd9f1eaa3;
    161: T0 = 32'hcd9fb7fb;
    162: T0 = 32'h4f163622;
    163: T0 = 32'h8377fcf2;
    164: T0 = 32'hc753f472;
    165: T0 = 32'hbf8d62d4;
    166: T0 = 32'hf5e1c59b;
    167: T0 = 32'ha4845b22;
    168: T0 = 32'h284e93b6;
    169: T0 = 32'h5f2d8e29;
    170: T0 = 32'h325a3f7a;
    171: T0 = 32'h9e45f195;
    172: T0 = 32'h665a81e7;
    173: T0 = 32'h7a5e5387;
    174: T0 = 32'ha5e9aa03;
    175: T0 = 32'h513c1499;
    176: T0 = 32'h6e827a66;
    177: T0 = 32'h95feae7c;
    178: T0 = 32'h658ba242;
    179: T0 = 32'hffec2dfe;
    180: T0 = 32'h492866b7;
    181: T0 = 32'h5308341c;
    182: T0 = 32'hefce3054;
    183: T0 = 32'h3db80e7f;
    184: T0 = 32'h93380515;
    185: T0 = 32'ha6e63902;
    186: T0 = 32'h81dd4fc0;
    187: T0 = 32'heb3f47f6;
    188: T0 = 32'h988f6690;
    189: T0 = 32'ha32f1720;
    190: T0 = 32'hd0ce559e;
    191: T0 = 32'hce414eaf;
    192: T0 = 32'hc1d76efd;
    193: T0 = 32'hc91dca12;
    194: T0 = 32'hf0ac0c8f;
    195: T0 = 32'hdc3db80a;
    196: T0 = 32'h72112505;
    197: T0 = 32'h1a8c7cc3;
    198: T0 = 32'haed78d2a;
    199: T0 = 32'hd61d48a7;
    200: T0 = 32'h71a0707b;
    201: T0 = 32'he9cb6756;
    202: T0 = 32'he0a7ba72;
    203: T0 = 32'h35cf2574;
    204: T0 = 32'ha6bd2ce6;
    205: T0 = 32'h936bbbca;
    206: T0 = 32'hc606bc30;
    207: T0 = 32'h62e276e8;
    208: T0 = 32'h717870b2;
    209: T0 = 32'he74275cb;
    210: T0 = 32'hcae6160e;
    211: T0 = 32'h834b20e8;
    212: T0 = 32'h6d7d6ea;
    213: T0 = 32'hce9d4bbf;
    214: T0 = 32'hf53843ff;
    215: T0 = 32'h30c0299a;
    216: T0 = 32'h182ea3da;
    217: T0 = 32'h898d83be;
    218: T0 = 32'h7b72077e;
    219: T0 = 32'h5d459019;
    220: T0 = 32'h4176512f;
    221: T0 = 32'h7a765263;
    222: T0 = 32'ha4e88283;
    223: T0 = 32'h53179cf5;
    224: T0 = 32'ha7869d79;
    225: T0 = 32'h3b4c9d13;
    226: T0 = 32'h10047d3f;
    227: T0 = 32'hc8ccb98a;
    228: T0 = 32'h93c014a;
    229: T0 = 32'h389f8c2;
    230: T0 = 32'h38af9f49;
    231: T0 = 32'hb275cc94;
    232: T0 = 32'h85f927eb;
    233: T0 = 32'h64c1a4d0;
    234: T0 = 32'hf984283b;
    235: T0 = 32'hc086ad22;
    236: T0 = 32'h9fea8888;
    237: T0 = 32'h6893d9d3;
    238: T0 = 32'h2d56ca74;
    239: T0 = 32'h94d8d0c9;
    240: T0 = 32'hea22c0cb;
    241: T0 = 32'heb8597eb;
    242: T0 = 32'h1701e2c5;
    243: T0 = 32'h71916ec1;
    244: T0 = 32'he744efad;
    245: T0 = 32'hd9f5c761;
    246: T0 = 32'h96040c8e;
    247: T0 = 32'h8e04730d;
    248: T0 = 32'h71ed9a28;
    249: T0 = 32'h5f5d1389;
    250: T0 = 32'h2613936d;
    251: T0 = 32'ha2b86895;
    252: T0 = 32'haaf4f777;
    253: T0 = 32'h9d4362c5;
    254: T0 = 32'h3bfd7b4e;
    255: T0 = 32'h29fb22d7;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[7:0];
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T6 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_25(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[7:0] io_weights
);

  reg [7:0] weightsReg;
  wire[7:0] T4;
  reg [7:0] T0;
  wire[7:0] T5;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T6;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 8'h0 : T0;
  always @(*) case (T5)
    0: T0 = 8'hf6;
    1: T0 = 8'hf5;
    2: T0 = 8'hf0;
    3: T0 = 8'hfc;
    4: T0 = 8'hf4;
    5: T0 = 8'h6;
    6: T0 = 8'he9;
    7: T0 = 8'h4;
    8: T0 = 8'hf;
    9: T0 = 8'h8;
    10: T0 = 8'hf1;
    11: T0 = 8'hd;
    12: T0 = 8'h6;
    13: T0 = 8'h10;
    14: T0 = 8'hf0;
    15: T0 = 8'hf4;
    16: T0 = 8'hff;
    17: T0 = 8'hf8;
    18: T0 = 8'he4;
    19: T0 = 8'hfb;
    20: T0 = 8'hf4;
    21: T0 = 8'h17;
    22: T0 = 8'h4;
    23: T0 = 8'h11;
    24: T0 = 8'h4;
    25: T0 = 8'h18;
    26: T0 = 8'he8;
    27: T0 = 8'ha;
    28: T0 = 8'hf;
    29: T0 = 8'h1;
    30: T0 = 8'h8;
    31: T0 = 8'hfc;
    32: T0 = 8'hf5;
    33: T0 = 8'hfd;
    34: T0 = 8'h1e;
    35: T0 = 8'h2;
    36: T0 = 8'h17;
    37: T0 = 8'hf3;
    38: T0 = 8'h5;
    39: T0 = 8'h2;
    40: T0 = 8'hf5;
    41: T0 = 8'h11;
    42: T0 = 8'hfe;
    43: T0 = 8'he;
    44: T0 = 8'ha;
    45: T0 = 8'hfa;
    46: T0 = 8'hec;
    47: T0 = 8'hfa;
    48: T0 = 8'h7;
    49: T0 = 8'hb;
    50: T0 = 8'hc;
    51: T0 = 8'hf2;
    52: T0 = 8'hf6;
    53: T0 = 8'hd;
    54: T0 = 8'hf5;
    55: T0 = 8'h4;
    56: T0 = 8'hee;
    57: T0 = 8'hf1;
    58: T0 = 8'h12;
    59: T0 = 8'hfa;
    60: T0 = 8'hfd;
    61: T0 = 8'h2;
    62: T0 = 8'hed;
    63: T0 = 8'h6;
    64: T0 = 8'hf0;
    65: T0 = 8'hf4;
    66: T0 = 8'hd;
    67: T0 = 8'hfa;
    68: T0 = 8'h0;
    69: T0 = 8'hfa;
    70: T0 = 8'hf4;
    71: T0 = 8'h1a;
    72: T0 = 8'h7;
    73: T0 = 8'hf;
    74: T0 = 8'he;
    75: T0 = 8'hff;
    76: T0 = 8'h0;
    77: T0 = 8'h0;
    78: T0 = 8'hf2;
    79: T0 = 8'h8;
    80: T0 = 8'h6;
    81: T0 = 8'hb;
    82: T0 = 8'hff;
    83: T0 = 8'hf5;
    84: T0 = 8'h9;
    85: T0 = 8'h6;
    86: T0 = 8'he5;
    87: T0 = 8'h6;
    88: T0 = 8'hef;
    89: T0 = 8'hc;
    90: T0 = 8'hf4;
    91: T0 = 8'h7;
    92: T0 = 8'hf;
    93: T0 = 8'h8;
    94: T0 = 8'h2;
    95: T0 = 8'h7;
    96: T0 = 8'hf9;
    97: T0 = 8'hec;
    98: T0 = 8'hf7;
    99: T0 = 8'hee;
    100: T0 = 8'hc;
    101: T0 = 8'hf4;
    102: T0 = 8'hff;
    103: T0 = 8'hf0;
    104: T0 = 8'h8;
    105: T0 = 8'h19;
    106: T0 = 8'hfb;
    107: T0 = 8'hfb;
    108: T0 = 8'hd;
    109: T0 = 8'hf8;
    110: T0 = 8'hed;
    111: T0 = 8'hfb;
    112: T0 = 8'hf2;
    113: T0 = 8'hf0;
    114: T0 = 8'h0;
    115: T0 = 8'hc;
    116: T0 = 8'hfd;
    117: T0 = 8'hf2;
    118: T0 = 8'hea;
    119: T0 = 8'hf3;
    120: T0 = 8'hf2;
    121: T0 = 8'hee;
    122: T0 = 8'h10;
    123: T0 = 8'h8;
    124: T0 = 8'h2;
    125: T0 = 8'ha;
    126: T0 = 8'h18;
    127: T0 = 8'hf2;
    128: T0 = 8'hef;
    129: T0 = 8'he;
    130: T0 = 8'he;
    131: T0 = 8'hf5;
    132: T0 = 8'hf7;
    133: T0 = 8'h12;
    134: T0 = 8'hf1;
    135: T0 = 8'hfe;
    136: T0 = 8'hfa;
    137: T0 = 8'heb;
    138: T0 = 8'h1c;
    139: T0 = 8'heb;
    140: T0 = 8'hd;
    141: T0 = 8'hf1;
    142: T0 = 8'hc;
    143: T0 = 8'h11;
    144: T0 = 8'hee;
    145: T0 = 8'hf2;
    146: T0 = 8'hf;
    147: T0 = 8'h7;
    148: T0 = 8'ha;
    149: T0 = 8'hf5;
    150: T0 = 8'hfe;
    151: T0 = 8'h9;
    152: T0 = 8'hec;
    153: T0 = 8'hf1;
    154: T0 = 8'h6;
    155: T0 = 8'h11;
    156: T0 = 8'h9;
    157: T0 = 8'hf5;
    158: T0 = 8'h1;
    159: T0 = 8'h0;
    160: T0 = 8'hed;
    161: T0 = 8'hf8;
    162: T0 = 8'hfe;
    163: T0 = 8'hfe;
    164: T0 = 8'hc;
    165: T0 = 8'h3;
    166: T0 = 8'he9;
    167: T0 = 8'hf0;
    168: T0 = 8'hf;
    169: T0 = 8'hf6;
    170: T0 = 8'h6;
    171: T0 = 8'h1;
    172: T0 = 8'hfd;
    173: T0 = 8'hf2;
    174: T0 = 8'h8;
    175: T0 = 8'he2;
    176: T0 = 8'hfc;
    177: T0 = 8'he2;
    178: T0 = 8'h0;
    179: T0 = 8'h1a;
    180: T0 = 8'hf2;
    181: T0 = 8'h3;
    182: T0 = 8'h8;
    183: T0 = 8'he;
    184: T0 = 8'h2;
    185: T0 = 8'h1;
    186: T0 = 8'hfa;
    187: T0 = 8'h6;
    188: T0 = 8'h14;
    189: T0 = 8'hfb;
    190: T0 = 8'hb;
    191: T0 = 8'he9;
    192: T0 = 8'hd7;
    193: T0 = 8'hc;
    194: T0 = 8'hd;
    195: T0 = 8'hf4;
    196: T0 = 8'h3;
    197: T0 = 8'hfe;
    198: T0 = 8'hf1;
    199: T0 = 8'ha;
    200: T0 = 8'hc;
    201: T0 = 8'h5;
    202: T0 = 8'h6;
    203: T0 = 8'hff;
    204: T0 = 8'hd;
    205: T0 = 8'hf6;
    206: T0 = 8'h7;
    207: T0 = 8'hf2;
    208: T0 = 8'h1;
    209: T0 = 8'hc;
    210: T0 = 8'hec;
    211: T0 = 8'h3;
    212: T0 = 8'h5;
    213: T0 = 8'hee;
    214: T0 = 8'hd;
    215: T0 = 8'hfc;
    216: T0 = 8'he;
    217: T0 = 8'h4;
    218: T0 = 8'h7;
    219: T0 = 8'hef;
    220: T0 = 8'h0;
    221: T0 = 8'he9;
    222: T0 = 8'he;
    223: T0 = 8'hf5;
    224: T0 = 8'hf0;
    225: T0 = 8'hc;
    226: T0 = 8'h5;
    227: T0 = 8'h10;
    228: T0 = 8'he5;
    229: T0 = 8'h10;
    230: T0 = 8'h9;
    231: T0 = 8'hfe;
    232: T0 = 8'ha;
    233: T0 = 8'h1b;
    234: T0 = 8'hf9;
    235: T0 = 8'h10;
    236: T0 = 8'h12;
    237: T0 = 8'hb;
    238: T0 = 8'h14;
    239: T0 = 8'hf4;
    240: T0 = 8'hed;
    241: T0 = 8'hfa;
    242: T0 = 8'hed;
    243: T0 = 8'h16;
    244: T0 = 8'hff;
    245: T0 = 8'hed;
    246: T0 = 8'h10;
    247: T0 = 8'h3;
    248: T0 = 8'hfc;
    249: T0 = 8'h10;
    250: T0 = 8'hf2;
    251: T0 = 8'hf3;
    252: T0 = 8'hf;
    253: T0 = 8'h15;
    254: T0 = 8'h3;
    255: T0 = 8'h4;
    default: begin
      T0 = 8'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[7:0];
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T6 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 8'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryStreamer_1(input clk, input reset,
    input  io_restart,
    output[15:0] io_weights_15,
    output[15:0] io_weights_14,
    output[15:0] io_weights_13,
    output[15:0] io_weights_12,
    output[15:0] io_weights_11,
    output[15:0] io_weights_10,
    output[15:0] io_weights_9,
    output[15:0] io_weights_8,
    output[15:0] io_weights_7,
    output[15:0] io_weights_6,
    output[15:0] io_weights_5,
    output[15:0] io_weights_4,
    output[15:0] io_weights_3,
    output[15:0] io_weights_2,
    output[15:0] io_weights_1,
    output[15:0] io_weights_0,
    output[7:0] io_bias
);

  wire[7:0] T18;
  wire[8:0] T0;
  wire[8:0] T1;
  wire[15:0] T2;
  wire[15:0] T3;
  wire[15:0] T4;
  wire[15:0] T5;
  wire[15:0] T6;
  wire[15:0] T7;
  wire[15:0] T8;
  wire[15:0] T9;
  wire[15:0] T10;
  wire[15:0] T11;
  wire[15:0] T12;
  wire[15:0] T13;
  wire[15:0] T14;
  wire[15:0] T15;
  wire[15:0] T16;
  wire[15:0] T17;
  wire MemoryUnit_io_restartOut;
  wire[31:0] MemoryUnit_io_weights;
  wire MemoryUnit_1_io_restartOut;
  wire[31:0] MemoryUnit_1_io_weights;
  wire MemoryUnit_2_io_restartOut;
  wire[31:0] MemoryUnit_2_io_weights;
  wire MemoryUnit_3_io_restartOut;
  wire[31:0] MemoryUnit_3_io_weights;
  wire MemoryUnit_4_io_restartOut;
  wire[31:0] MemoryUnit_4_io_weights;
  wire MemoryUnit_5_io_restartOut;
  wire[31:0] MemoryUnit_5_io_weights;
  wire MemoryUnit_6_io_restartOut;
  wire[31:0] MemoryUnit_6_io_weights;
  wire[31:0] MemoryUnit_7_io_weights;
  wire[7:0] biasMemoryUnit_io_weights;


  assign io_bias = T18;
  assign T18 = T0[7:0];
  assign T0 = T1;
  assign T1 = {1'h0, biasMemoryUnit_io_weights};
  assign io_weights_0 = T2;
  assign T2 = MemoryUnit_io_weights[15:0];
  assign io_weights_1 = T3;
  assign T3 = MemoryUnit_io_weights[31:16];
  assign io_weights_2 = T4;
  assign T4 = MemoryUnit_1_io_weights[15:0];
  assign io_weights_3 = T5;
  assign T5 = MemoryUnit_1_io_weights[31:16];
  assign io_weights_4 = T6;
  assign T6 = MemoryUnit_2_io_weights[15:0];
  assign io_weights_5 = T7;
  assign T7 = MemoryUnit_2_io_weights[31:16];
  assign io_weights_6 = T8;
  assign T8 = MemoryUnit_3_io_weights[15:0];
  assign io_weights_7 = T9;
  assign T9 = MemoryUnit_3_io_weights[31:16];
  assign io_weights_8 = T10;
  assign T10 = MemoryUnit_4_io_weights[15:0];
  assign io_weights_9 = T11;
  assign T11 = MemoryUnit_4_io_weights[31:16];
  assign io_weights_10 = T12;
  assign T12 = MemoryUnit_5_io_weights[15:0];
  assign io_weights_11 = T13;
  assign T13 = MemoryUnit_5_io_weights[31:16];
  assign io_weights_12 = T14;
  assign T14 = MemoryUnit_6_io_weights[15:0];
  assign io_weights_13 = T15;
  assign T15 = MemoryUnit_6_io_weights[31:16];
  assign io_weights_14 = T16;
  assign T16 = MemoryUnit_7_io_weights[15:0];
  assign io_weights_15 = T17;
  assign T17 = MemoryUnit_7_io_weights[31:16];
  MemoryUnit_17 MemoryUnit(.clk(clk), .reset(reset),
       .io_restartIn( io_restart ),
       .io_restartOut( MemoryUnit_io_restartOut ),
       .io_weights( MemoryUnit_io_weights )
  );
  MemoryUnit_18 MemoryUnit_1(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_io_restartOut ),
       .io_restartOut( MemoryUnit_1_io_restartOut ),
       .io_weights( MemoryUnit_1_io_weights )
  );
  MemoryUnit_19 MemoryUnit_2(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_1_io_restartOut ),
       .io_restartOut( MemoryUnit_2_io_restartOut ),
       .io_weights( MemoryUnit_2_io_weights )
  );
  MemoryUnit_20 MemoryUnit_3(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_2_io_restartOut ),
       .io_restartOut( MemoryUnit_3_io_restartOut ),
       .io_weights( MemoryUnit_3_io_weights )
  );
  MemoryUnit_21 MemoryUnit_4(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_3_io_restartOut ),
       .io_restartOut( MemoryUnit_4_io_restartOut ),
       .io_weights( MemoryUnit_4_io_weights )
  );
  MemoryUnit_22 MemoryUnit_5(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_4_io_restartOut ),
       .io_restartOut( MemoryUnit_5_io_restartOut ),
       .io_weights( MemoryUnit_5_io_weights )
  );
  MemoryUnit_23 MemoryUnit_6(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_5_io_restartOut ),
       .io_restartOut( MemoryUnit_6_io_restartOut ),
       .io_weights( MemoryUnit_6_io_weights )
  );
  MemoryUnit_24 MemoryUnit_7(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_6_io_restartOut ),
       //.io_restartOut(  )
       .io_weights( MemoryUnit_7_io_weights )
  );
  MemoryUnit_25 biasMemoryUnit(.clk(clk), .reset(reset),
       .io_restartIn( io_restart ),
       //.io_restartOut(  )
       .io_weights( biasMemoryUnit_io_weights )
  );
endmodule

module Warp_1(input clk, input reset,
    input [15:0] io_xIn_2,
    input [15:0] io_xIn_1,
    input [15:0] io_xIn_0,
    input  io_start,
    output io_ready,
    output io_startOut,
    output io_xOut_2,
    output io_xOut_1,
    output io_xOut_0,
    output io_xOutValid,
    input  io_pipeReady,
    output io_done
);

  wire[9:0] T189;
  wire[10:0] T0;
  wire[10:0] T1;
  wire[9:0] T190;
  wire[10:0] T2;
  wire[10:0] T3;
  wire[9:0] T191;
  wire[10:0] T4;
  wire[10:0] T5;
  wire[9:0] T192;
  wire[10:0] T6;
  wire[10:0] T7;
  wire[9:0] T193;
  wire[10:0] T8;
  wire[10:0] T9;
  wire[9:0] T194;
  wire[10:0] T10;
  wire[10:0] T11;
  wire[9:0] T195;
  wire[10:0] T12;
  wire[10:0] T13;
  wire[9:0] T196;
  wire[10:0] T14;
  wire[10:0] T15;
  wire[9:0] T197;
  wire[10:0] T16;
  wire[10:0] T17;
  wire[9:0] T198;
  wire[10:0] T18;
  wire[10:0] T19;
  wire[9:0] T199;
  wire[10:0] T20;
  wire[10:0] T21;
  wire[9:0] T200;
  wire[10:0] T22;
  wire[10:0] T23;
  wire[9:0] T201;
  wire[10:0] T24;
  wire[10:0] T25;
  wire[9:0] T202;
  wire[10:0] T26;
  wire[10:0] T27;
  wire[9:0] T203;
  wire[10:0] T28;
  wire[10:0] T29;
  wire[9:0] T204;
  wire[10:0] T30;
  wire[10:0] T31;
  wire[9:0] T205;
  wire[10:0] T32;
  wire[10:0] T33;
  wire[9:0] T206;
  wire[10:0] T34;
  wire[10:0] T35;
  wire[9:0] T207;
  wire[10:0] T36;
  wire[10:0] T37;
  wire[9:0] T208;
  wire[10:0] T38;
  wire[10:0] T39;
  wire[9:0] T209;
  wire[10:0] T40;
  wire[10:0] T41;
  wire[9:0] T210;
  wire[10:0] T42;
  wire[10:0] T43;
  wire[9:0] T211;
  wire[10:0] T44;
  wire[10:0] T45;
  wire[9:0] T212;
  wire[10:0] T46;
  wire[10:0] T47;
  wire[9:0] T213;
  wire[10:0] T48;
  wire[10:0] T49;
  wire[9:0] T214;
  wire[10:0] T50;
  wire[10:0] T51;
  wire[9:0] T215;
  wire[10:0] T52;
  wire[10:0] T53;
  wire[9:0] T216;
  wire[10:0] T54;
  wire[10:0] T55;
  wire[9:0] T217;
  wire[10:0] T56;
  wire[10:0] T57;
  wire[9:0] T218;
  wire[10:0] T58;
  wire[10:0] T59;
  wire[9:0] T219;
  wire[10:0] T60;
  wire[10:0] T61;
  wire[9:0] T220;
  wire[10:0] T62;
  wire[10:0] T63;
  wire[9:0] T221;
  wire[10:0] T64;
  wire[10:0] T65;
  wire[9:0] T222;
  wire[10:0] T66;
  wire[10:0] T67;
  wire[9:0] T223;
  wire[10:0] T68;
  wire[10:0] T69;
  wire[9:0] T224;
  wire[10:0] T70;
  wire[10:0] T71;
  wire[9:0] T225;
  wire[10:0] T72;
  wire[10:0] T73;
  wire[9:0] T226;
  wire[10:0] T74;
  wire[10:0] T75;
  wire[9:0] T227;
  wire[10:0] T76;
  wire[10:0] T77;
  wire[9:0] T228;
  wire[10:0] T78;
  wire[10:0] T79;
  wire[9:0] T229;
  wire[10:0] T80;
  wire[10:0] T81;
  wire[9:0] T230;
  wire[10:0] T82;
  wire[10:0] T83;
  wire[9:0] T231;
  wire[10:0] T84;
  wire[10:0] T85;
  wire[9:0] T232;
  wire[10:0] T86;
  wire[10:0] T87;
  wire[9:0] T233;
  wire[10:0] T88;
  wire[10:0] T89;
  wire[9:0] T234;
  wire[10:0] T90;
  wire[10:0] T91;
  wire[9:0] T235;
  wire[10:0] T92;
  wire[10:0] T93;
  wire[9:0] T236;
  wire[10:0] T94;
  wire[10:0] T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire[3:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire[3:0] T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire[3:0] T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire Activation_io_out_15;
  wire Activation_io_out_14;
  wire Activation_io_out_13;
  wire Activation_io_out_12;
  wire Activation_io_out_11;
  wire Activation_io_out_10;
  wire Activation_io_out_9;
  wire Activation_io_out_8;
  wire Activation_io_out_7;
  wire Activation_io_out_6;
  wire Activation_io_out_5;
  wire Activation_io_out_4;
  wire Activation_io_out_3;
  wire Activation_io_out_2;
  wire Activation_io_out_1;
  wire Activation_io_out_0;
  wire Activation_1_io_out_15;
  wire Activation_1_io_out_14;
  wire Activation_1_io_out_13;
  wire Activation_1_io_out_12;
  wire Activation_1_io_out_11;
  wire Activation_1_io_out_10;
  wire Activation_1_io_out_9;
  wire Activation_1_io_out_8;
  wire Activation_1_io_out_7;
  wire Activation_1_io_out_6;
  wire Activation_1_io_out_5;
  wire Activation_1_io_out_4;
  wire Activation_1_io_out_3;
  wire Activation_1_io_out_2;
  wire Activation_1_io_out_1;
  wire Activation_1_io_out_0;
  wire Activation_2_io_out_15;
  wire Activation_2_io_out_14;
  wire Activation_2_io_out_13;
  wire Activation_2_io_out_12;
  wire Activation_2_io_out_11;
  wire Activation_2_io_out_10;
  wire Activation_2_io_out_9;
  wire Activation_2_io_out_8;
  wire Activation_2_io_out_7;
  wire Activation_2_io_out_6;
  wire Activation_2_io_out_5;
  wire Activation_2_io_out_4;
  wire Activation_2_io_out_3;
  wire Activation_2_io_out_2;
  wire Activation_2_io_out_1;
  wire Activation_2_io_out_0;
  wire control_io_ready;
  wire control_io_valid;
  wire control_io_done;
  wire[3:0] control_io_selectX;
  wire control_io_memoryRestart;
  wire control_io_chainRestart;
  wire[9:0] Chain_io_ys_15;
  wire[9:0] Chain_io_ys_14;
  wire[9:0] Chain_io_ys_13;
  wire[9:0] Chain_io_ys_12;
  wire[9:0] Chain_io_ys_11;
  wire[9:0] Chain_io_ys_10;
  wire[9:0] Chain_io_ys_9;
  wire[9:0] Chain_io_ys_8;
  wire[9:0] Chain_io_ys_7;
  wire[9:0] Chain_io_ys_6;
  wire[9:0] Chain_io_ys_5;
  wire[9:0] Chain_io_ys_4;
  wire[9:0] Chain_io_ys_3;
  wire[9:0] Chain_io_ys_2;
  wire[9:0] Chain_io_ys_1;
  wire[9:0] Chain_io_ys_0;
  wire[9:0] Chain_1_io_ys_15;
  wire[9:0] Chain_1_io_ys_14;
  wire[9:0] Chain_1_io_ys_13;
  wire[9:0] Chain_1_io_ys_12;
  wire[9:0] Chain_1_io_ys_11;
  wire[9:0] Chain_1_io_ys_10;
  wire[9:0] Chain_1_io_ys_9;
  wire[9:0] Chain_1_io_ys_8;
  wire[9:0] Chain_1_io_ys_7;
  wire[9:0] Chain_1_io_ys_6;
  wire[9:0] Chain_1_io_ys_5;
  wire[9:0] Chain_1_io_ys_4;
  wire[9:0] Chain_1_io_ys_3;
  wire[9:0] Chain_1_io_ys_2;
  wire[9:0] Chain_1_io_ys_1;
  wire[9:0] Chain_1_io_ys_0;
  wire[9:0] Chain_2_io_ys_15;
  wire[9:0] Chain_2_io_ys_14;
  wire[9:0] Chain_2_io_ys_13;
  wire[9:0] Chain_2_io_ys_12;
  wire[9:0] Chain_2_io_ys_11;
  wire[9:0] Chain_2_io_ys_10;
  wire[9:0] Chain_2_io_ys_9;
  wire[9:0] Chain_2_io_ys_8;
  wire[9:0] Chain_2_io_ys_7;
  wire[9:0] Chain_2_io_ys_6;
  wire[9:0] Chain_2_io_ys_5;
  wire[9:0] Chain_2_io_ys_4;
  wire[9:0] Chain_2_io_ys_3;
  wire[9:0] Chain_2_io_ys_2;
  wire[9:0] Chain_2_io_ys_1;
  wire[9:0] Chain_2_io_ys_0;
  wire[15:0] memoryStreamer_io_weights_15;
  wire[15:0] memoryStreamer_io_weights_14;
  wire[15:0] memoryStreamer_io_weights_13;
  wire[15:0] memoryStreamer_io_weights_12;
  wire[15:0] memoryStreamer_io_weights_11;
  wire[15:0] memoryStreamer_io_weights_10;
  wire[15:0] memoryStreamer_io_weights_9;
  wire[15:0] memoryStreamer_io_weights_8;
  wire[15:0] memoryStreamer_io_weights_7;
  wire[15:0] memoryStreamer_io_weights_6;
  wire[15:0] memoryStreamer_io_weights_5;
  wire[15:0] memoryStreamer_io_weights_4;
  wire[15:0] memoryStreamer_io_weights_3;
  wire[15:0] memoryStreamer_io_weights_2;
  wire[15:0] memoryStreamer_io_weights_1;
  wire[15:0] memoryStreamer_io_weights_0;
  wire[7:0] memoryStreamer_io_bias;


  assign T189 = T0[9:0];
  assign T0 = T1;
  assign T1 = {1'h0, Chain_2_io_ys_0};
  assign T190 = T2[9:0];
  assign T2 = T3;
  assign T3 = {1'h0, Chain_2_io_ys_1};
  assign T191 = T4[9:0];
  assign T4 = T5;
  assign T5 = {1'h0, Chain_2_io_ys_2};
  assign T192 = T6[9:0];
  assign T6 = T7;
  assign T7 = {1'h0, Chain_2_io_ys_3};
  assign T193 = T8[9:0];
  assign T8 = T9;
  assign T9 = {1'h0, Chain_2_io_ys_4};
  assign T194 = T10[9:0];
  assign T10 = T11;
  assign T11 = {1'h0, Chain_2_io_ys_5};
  assign T195 = T12[9:0];
  assign T12 = T13;
  assign T13 = {1'h0, Chain_2_io_ys_6};
  assign T196 = T14[9:0];
  assign T14 = T15;
  assign T15 = {1'h0, Chain_2_io_ys_7};
  assign T197 = T16[9:0];
  assign T16 = T17;
  assign T17 = {1'h0, Chain_2_io_ys_8};
  assign T198 = T18[9:0];
  assign T18 = T19;
  assign T19 = {1'h0, Chain_2_io_ys_9};
  assign T199 = T20[9:0];
  assign T20 = T21;
  assign T21 = {1'h0, Chain_2_io_ys_10};
  assign T200 = T22[9:0];
  assign T22 = T23;
  assign T23 = {1'h0, Chain_2_io_ys_11};
  assign T201 = T24[9:0];
  assign T24 = T25;
  assign T25 = {1'h0, Chain_2_io_ys_12};
  assign T202 = T26[9:0];
  assign T26 = T27;
  assign T27 = {1'h0, Chain_2_io_ys_13};
  assign T203 = T28[9:0];
  assign T28 = T29;
  assign T29 = {1'h0, Chain_2_io_ys_14};
  assign T204 = T30[9:0];
  assign T30 = T31;
  assign T31 = {1'h0, Chain_2_io_ys_15};
  assign T205 = T32[9:0];
  assign T32 = T33;
  assign T33 = {1'h0, Chain_1_io_ys_0};
  assign T206 = T34[9:0];
  assign T34 = T35;
  assign T35 = {1'h0, Chain_1_io_ys_1};
  assign T207 = T36[9:0];
  assign T36 = T37;
  assign T37 = {1'h0, Chain_1_io_ys_2};
  assign T208 = T38[9:0];
  assign T38 = T39;
  assign T39 = {1'h0, Chain_1_io_ys_3};
  assign T209 = T40[9:0];
  assign T40 = T41;
  assign T41 = {1'h0, Chain_1_io_ys_4};
  assign T210 = T42[9:0];
  assign T42 = T43;
  assign T43 = {1'h0, Chain_1_io_ys_5};
  assign T211 = T44[9:0];
  assign T44 = T45;
  assign T45 = {1'h0, Chain_1_io_ys_6};
  assign T212 = T46[9:0];
  assign T46 = T47;
  assign T47 = {1'h0, Chain_1_io_ys_7};
  assign T213 = T48[9:0];
  assign T48 = T49;
  assign T49 = {1'h0, Chain_1_io_ys_8};
  assign T214 = T50[9:0];
  assign T50 = T51;
  assign T51 = {1'h0, Chain_1_io_ys_9};
  assign T215 = T52[9:0];
  assign T52 = T53;
  assign T53 = {1'h0, Chain_1_io_ys_10};
  assign T216 = T54[9:0];
  assign T54 = T55;
  assign T55 = {1'h0, Chain_1_io_ys_11};
  assign T217 = T56[9:0];
  assign T56 = T57;
  assign T57 = {1'h0, Chain_1_io_ys_12};
  assign T218 = T58[9:0];
  assign T58 = T59;
  assign T59 = {1'h0, Chain_1_io_ys_13};
  assign T219 = T60[9:0];
  assign T60 = T61;
  assign T61 = {1'h0, Chain_1_io_ys_14};
  assign T220 = T62[9:0];
  assign T62 = T63;
  assign T63 = {1'h0, Chain_1_io_ys_15};
  assign T221 = T64[9:0];
  assign T64 = T65;
  assign T65 = {1'h0, Chain_io_ys_0};
  assign T222 = T66[9:0];
  assign T66 = T67;
  assign T67 = {1'h0, Chain_io_ys_1};
  assign T223 = T68[9:0];
  assign T68 = T69;
  assign T69 = {1'h0, Chain_io_ys_2};
  assign T224 = T70[9:0];
  assign T70 = T71;
  assign T71 = {1'h0, Chain_io_ys_3};
  assign T225 = T72[9:0];
  assign T72 = T73;
  assign T73 = {1'h0, Chain_io_ys_4};
  assign T226 = T74[9:0];
  assign T74 = T75;
  assign T75 = {1'h0, Chain_io_ys_5};
  assign T227 = T76[9:0];
  assign T76 = T77;
  assign T77 = {1'h0, Chain_io_ys_6};
  assign T228 = T78[9:0];
  assign T78 = T79;
  assign T79 = {1'h0, Chain_io_ys_7};
  assign T229 = T80[9:0];
  assign T80 = T81;
  assign T81 = {1'h0, Chain_io_ys_8};
  assign T230 = T82[9:0];
  assign T82 = T83;
  assign T83 = {1'h0, Chain_io_ys_9};
  assign T231 = T84[9:0];
  assign T84 = T85;
  assign T85 = {1'h0, Chain_io_ys_10};
  assign T232 = T86[9:0];
  assign T86 = T87;
  assign T87 = {1'h0, Chain_io_ys_11};
  assign T233 = T88[9:0];
  assign T88 = T89;
  assign T89 = {1'h0, Chain_io_ys_12};
  assign T234 = T90[9:0];
  assign T90 = T91;
  assign T91 = {1'h0, Chain_io_ys_13};
  assign T235 = T92[9:0];
  assign T92 = T93;
  assign T93 = {1'h0, Chain_io_ys_14};
  assign T236 = T94[9:0];
  assign T94 = T95;
  assign T95 = {1'h0, Chain_io_ys_15};
  assign io_done = control_io_done;
  assign io_xOutValid = control_io_valid;
  assign io_xOut_0 = T96;
  assign T96 = T126 ? T112 : T97;
  assign T97 = T111 ? T105 : T98;
  assign T98 = T104 ? T102 : T99;
  assign T99 = T100 ? Activation_io_out_1 : Activation_io_out_0;
  assign T100 = T101[0];
  assign T101 = control_io_selectX;
  assign T102 = T103 ? Activation_io_out_3 : Activation_io_out_2;
  assign T103 = T101[0];
  assign T104 = T101[1];
  assign T105 = T110 ? T108 : T106;
  assign T106 = T107 ? Activation_io_out_5 : Activation_io_out_4;
  assign T107 = T101[0];
  assign T108 = T109 ? Activation_io_out_7 : Activation_io_out_6;
  assign T109 = T101[0];
  assign T110 = T101[1];
  assign T111 = T101[2];
  assign T112 = T125 ? T119 : T113;
  assign T113 = T118 ? T116 : T114;
  assign T114 = T115 ? Activation_io_out_9 : Activation_io_out_8;
  assign T115 = T101[0];
  assign T116 = T117 ? Activation_io_out_11 : Activation_io_out_10;
  assign T117 = T101[0];
  assign T118 = T101[1];
  assign T119 = T124 ? T122 : T120;
  assign T120 = T121 ? Activation_io_out_13 : Activation_io_out_12;
  assign T121 = T101[0];
  assign T122 = T123 ? Activation_io_out_15 : Activation_io_out_14;
  assign T123 = T101[0];
  assign T124 = T101[1];
  assign T125 = T101[2];
  assign T126 = T101[3];
  assign io_xOut_1 = T127;
  assign T127 = T157 ? T143 : T128;
  assign T128 = T142 ? T136 : T129;
  assign T129 = T135 ? T133 : T130;
  assign T130 = T131 ? Activation_1_io_out_1 : Activation_1_io_out_0;
  assign T131 = T132[0];
  assign T132 = control_io_selectX;
  assign T133 = T134 ? Activation_1_io_out_3 : Activation_1_io_out_2;
  assign T134 = T132[0];
  assign T135 = T132[1];
  assign T136 = T141 ? T139 : T137;
  assign T137 = T138 ? Activation_1_io_out_5 : Activation_1_io_out_4;
  assign T138 = T132[0];
  assign T139 = T140 ? Activation_1_io_out_7 : Activation_1_io_out_6;
  assign T140 = T132[0];
  assign T141 = T132[1];
  assign T142 = T132[2];
  assign T143 = T156 ? T150 : T144;
  assign T144 = T149 ? T147 : T145;
  assign T145 = T146 ? Activation_1_io_out_9 : Activation_1_io_out_8;
  assign T146 = T132[0];
  assign T147 = T148 ? Activation_1_io_out_11 : Activation_1_io_out_10;
  assign T148 = T132[0];
  assign T149 = T132[1];
  assign T150 = T155 ? T153 : T151;
  assign T151 = T152 ? Activation_1_io_out_13 : Activation_1_io_out_12;
  assign T152 = T132[0];
  assign T153 = T154 ? Activation_1_io_out_15 : Activation_1_io_out_14;
  assign T154 = T132[0];
  assign T155 = T132[1];
  assign T156 = T132[2];
  assign T157 = T132[3];
  assign io_xOut_2 = T158;
  assign T158 = T188 ? T174 : T159;
  assign T159 = T173 ? T167 : T160;
  assign T160 = T166 ? T164 : T161;
  assign T161 = T162 ? Activation_2_io_out_1 : Activation_2_io_out_0;
  assign T162 = T163[0];
  assign T163 = control_io_selectX;
  assign T164 = T165 ? Activation_2_io_out_3 : Activation_2_io_out_2;
  assign T165 = T163[0];
  assign T166 = T163[1];
  assign T167 = T172 ? T170 : T168;
  assign T168 = T169 ? Activation_2_io_out_5 : Activation_2_io_out_4;
  assign T169 = T163[0];
  assign T170 = T171 ? Activation_2_io_out_7 : Activation_2_io_out_6;
  assign T171 = T163[0];
  assign T172 = T163[1];
  assign T173 = T163[2];
  assign T174 = T187 ? T181 : T175;
  assign T175 = T180 ? T178 : T176;
  assign T176 = T177 ? Activation_2_io_out_9 : Activation_2_io_out_8;
  assign T177 = T163[0];
  assign T178 = T179 ? Activation_2_io_out_11 : Activation_2_io_out_10;
  assign T179 = T163[0];
  assign T180 = T163[1];
  assign T181 = T186 ? T184 : T182;
  assign T182 = T183 ? Activation_2_io_out_13 : Activation_2_io_out_12;
  assign T183 = T163[0];
  assign T184 = T185 ? Activation_2_io_out_15 : Activation_2_io_out_14;
  assign T185 = T163[0];
  assign T186 = T163[1];
  assign T187 = T163[2];
  assign T188 = T163[3];
  assign io_startOut = io_start;
  assign io_ready = control_io_ready;
  WarpControl_1 control(.clk(clk), .reset(reset),
       .io_ready( control_io_ready ),
       .io_start( io_start ),
       .io_nextReady( io_pipeReady ),
       .io_valid( control_io_valid ),
       .io_done( control_io_done ),
       .io_selectX( control_io_selectX ),
       .io_memoryRestart( control_io_memoryRestart ),
       .io_chainRestart( control_io_chainRestart )
  );
  Chain_1 Chain(.clk(clk), .reset(reset),
       .io_weights_15( memoryStreamer_io_weights_15 ),
       .io_weights_14( memoryStreamer_io_weights_14 ),
       .io_weights_13( memoryStreamer_io_weights_13 ),
       .io_weights_12( memoryStreamer_io_weights_12 ),
       .io_weights_11( memoryStreamer_io_weights_11 ),
       .io_weights_10( memoryStreamer_io_weights_10 ),
       .io_weights_9( memoryStreamer_io_weights_9 ),
       .io_weights_8( memoryStreamer_io_weights_8 ),
       .io_weights_7( memoryStreamer_io_weights_7 ),
       .io_weights_6( memoryStreamer_io_weights_6 ),
       .io_weights_5( memoryStreamer_io_weights_5 ),
       .io_weights_4( memoryStreamer_io_weights_4 ),
       .io_weights_3( memoryStreamer_io_weights_3 ),
       .io_weights_2( memoryStreamer_io_weights_2 ),
       .io_weights_1( memoryStreamer_io_weights_1 ),
       .io_weights_0( memoryStreamer_io_weights_0 ),
       .io_bias( memoryStreamer_io_bias ),
       .io_restartIn( control_io_chainRestart ),
       .io_xs( io_xIn_0 ),
       .io_ys_15( Chain_io_ys_15 ),
       .io_ys_14( Chain_io_ys_14 ),
       .io_ys_13( Chain_io_ys_13 ),
       .io_ys_12( Chain_io_ys_12 ),
       .io_ys_11( Chain_io_ys_11 ),
       .io_ys_10( Chain_io_ys_10 ),
       .io_ys_9( Chain_io_ys_9 ),
       .io_ys_8( Chain_io_ys_8 ),
       .io_ys_7( Chain_io_ys_7 ),
       .io_ys_6( Chain_io_ys_6 ),
       .io_ys_5( Chain_io_ys_5 ),
       .io_ys_4( Chain_io_ys_4 ),
       .io_ys_3( Chain_io_ys_3 ),
       .io_ys_2( Chain_io_ys_2 ),
       .io_ys_1( Chain_io_ys_1 ),
       .io_ys_0( Chain_io_ys_0 )
  );
  Chain_1 Chain_1(.clk(clk), .reset(reset),
       .io_weights_15( memoryStreamer_io_weights_15 ),
       .io_weights_14( memoryStreamer_io_weights_14 ),
       .io_weights_13( memoryStreamer_io_weights_13 ),
       .io_weights_12( memoryStreamer_io_weights_12 ),
       .io_weights_11( memoryStreamer_io_weights_11 ),
       .io_weights_10( memoryStreamer_io_weights_10 ),
       .io_weights_9( memoryStreamer_io_weights_9 ),
       .io_weights_8( memoryStreamer_io_weights_8 ),
       .io_weights_7( memoryStreamer_io_weights_7 ),
       .io_weights_6( memoryStreamer_io_weights_6 ),
       .io_weights_5( memoryStreamer_io_weights_5 ),
       .io_weights_4( memoryStreamer_io_weights_4 ),
       .io_weights_3( memoryStreamer_io_weights_3 ),
       .io_weights_2( memoryStreamer_io_weights_2 ),
       .io_weights_1( memoryStreamer_io_weights_1 ),
       .io_weights_0( memoryStreamer_io_weights_0 ),
       .io_bias( memoryStreamer_io_bias ),
       .io_restartIn( control_io_chainRestart ),
       .io_xs( io_xIn_1 ),
       .io_ys_15( Chain_1_io_ys_15 ),
       .io_ys_14( Chain_1_io_ys_14 ),
       .io_ys_13( Chain_1_io_ys_13 ),
       .io_ys_12( Chain_1_io_ys_12 ),
       .io_ys_11( Chain_1_io_ys_11 ),
       .io_ys_10( Chain_1_io_ys_10 ),
       .io_ys_9( Chain_1_io_ys_9 ),
       .io_ys_8( Chain_1_io_ys_8 ),
       .io_ys_7( Chain_1_io_ys_7 ),
       .io_ys_6( Chain_1_io_ys_6 ),
       .io_ys_5( Chain_1_io_ys_5 ),
       .io_ys_4( Chain_1_io_ys_4 ),
       .io_ys_3( Chain_1_io_ys_3 ),
       .io_ys_2( Chain_1_io_ys_2 ),
       .io_ys_1( Chain_1_io_ys_1 ),
       .io_ys_0( Chain_1_io_ys_0 )
  );
  Chain_1 Chain_2(.clk(clk), .reset(reset),
       .io_weights_15( memoryStreamer_io_weights_15 ),
       .io_weights_14( memoryStreamer_io_weights_14 ),
       .io_weights_13( memoryStreamer_io_weights_13 ),
       .io_weights_12( memoryStreamer_io_weights_12 ),
       .io_weights_11( memoryStreamer_io_weights_11 ),
       .io_weights_10( memoryStreamer_io_weights_10 ),
       .io_weights_9( memoryStreamer_io_weights_9 ),
       .io_weights_8( memoryStreamer_io_weights_8 ),
       .io_weights_7( memoryStreamer_io_weights_7 ),
       .io_weights_6( memoryStreamer_io_weights_6 ),
       .io_weights_5( memoryStreamer_io_weights_5 ),
       .io_weights_4( memoryStreamer_io_weights_4 ),
       .io_weights_3( memoryStreamer_io_weights_3 ),
       .io_weights_2( memoryStreamer_io_weights_2 ),
       .io_weights_1( memoryStreamer_io_weights_1 ),
       .io_weights_0( memoryStreamer_io_weights_0 ),
       .io_bias( memoryStreamer_io_bias ),
       .io_restartIn( control_io_chainRestart ),
       .io_xs( io_xIn_2 ),
       .io_ys_15( Chain_2_io_ys_15 ),
       .io_ys_14( Chain_2_io_ys_14 ),
       .io_ys_13( Chain_2_io_ys_13 ),
       .io_ys_12( Chain_2_io_ys_12 ),
       .io_ys_11( Chain_2_io_ys_11 ),
       .io_ys_10( Chain_2_io_ys_10 ),
       .io_ys_9( Chain_2_io_ys_9 ),
       .io_ys_8( Chain_2_io_ys_8 ),
       .io_ys_7( Chain_2_io_ys_7 ),
       .io_ys_6( Chain_2_io_ys_6 ),
       .io_ys_5( Chain_2_io_ys_5 ),
       .io_ys_4( Chain_2_io_ys_4 ),
       .io_ys_3( Chain_2_io_ys_3 ),
       .io_ys_2( Chain_2_io_ys_2 ),
       .io_ys_1( Chain_2_io_ys_1 ),
       .io_ys_0( Chain_2_io_ys_0 )
  );
  Activation_1 Activation(
       .io_in_15( T236 ),
       .io_in_14( T235 ),
       .io_in_13( T234 ),
       .io_in_12( T233 ),
       .io_in_11( T232 ),
       .io_in_10( T231 ),
       .io_in_9( T230 ),
       .io_in_8( T229 ),
       .io_in_7( T228 ),
       .io_in_6( T227 ),
       .io_in_5( T226 ),
       .io_in_4( T225 ),
       .io_in_3( T224 ),
       .io_in_2( T223 ),
       .io_in_1( T222 ),
       .io_in_0( T221 ),
       .io_out_15( Activation_io_out_15 ),
       .io_out_14( Activation_io_out_14 ),
       .io_out_13( Activation_io_out_13 ),
       .io_out_12( Activation_io_out_12 ),
       .io_out_11( Activation_io_out_11 ),
       .io_out_10( Activation_io_out_10 ),
       .io_out_9( Activation_io_out_9 ),
       .io_out_8( Activation_io_out_8 ),
       .io_out_7( Activation_io_out_7 ),
       .io_out_6( Activation_io_out_6 ),
       .io_out_5( Activation_io_out_5 ),
       .io_out_4( Activation_io_out_4 ),
       .io_out_3( Activation_io_out_3 ),
       .io_out_2( Activation_io_out_2 ),
       .io_out_1( Activation_io_out_1 ),
       .io_out_0( Activation_io_out_0 )
  );
  Activation_1 Activation_1(
       .io_in_15( T220 ),
       .io_in_14( T219 ),
       .io_in_13( T218 ),
       .io_in_12( T217 ),
       .io_in_11( T216 ),
       .io_in_10( T215 ),
       .io_in_9( T214 ),
       .io_in_8( T213 ),
       .io_in_7( T212 ),
       .io_in_6( T211 ),
       .io_in_5( T210 ),
       .io_in_4( T209 ),
       .io_in_3( T208 ),
       .io_in_2( T207 ),
       .io_in_1( T206 ),
       .io_in_0( T205 ),
       .io_out_15( Activation_1_io_out_15 ),
       .io_out_14( Activation_1_io_out_14 ),
       .io_out_13( Activation_1_io_out_13 ),
       .io_out_12( Activation_1_io_out_12 ),
       .io_out_11( Activation_1_io_out_11 ),
       .io_out_10( Activation_1_io_out_10 ),
       .io_out_9( Activation_1_io_out_9 ),
       .io_out_8( Activation_1_io_out_8 ),
       .io_out_7( Activation_1_io_out_7 ),
       .io_out_6( Activation_1_io_out_6 ),
       .io_out_5( Activation_1_io_out_5 ),
       .io_out_4( Activation_1_io_out_4 ),
       .io_out_3( Activation_1_io_out_3 ),
       .io_out_2( Activation_1_io_out_2 ),
       .io_out_1( Activation_1_io_out_1 ),
       .io_out_0( Activation_1_io_out_0 )
  );
  Activation_1 Activation_2(
       .io_in_15( T204 ),
       .io_in_14( T203 ),
       .io_in_13( T202 ),
       .io_in_12( T201 ),
       .io_in_11( T200 ),
       .io_in_10( T199 ),
       .io_in_9( T198 ),
       .io_in_8( T197 ),
       .io_in_7( T196 ),
       .io_in_6( T195 ),
       .io_in_5( T194 ),
       .io_in_4( T193 ),
       .io_in_3( T192 ),
       .io_in_2( T191 ),
       .io_in_1( T190 ),
       .io_in_0( T189 ),
       .io_out_15( Activation_2_io_out_15 ),
       .io_out_14( Activation_2_io_out_14 ),
       .io_out_13( Activation_2_io_out_13 ),
       .io_out_12( Activation_2_io_out_12 ),
       .io_out_11( Activation_2_io_out_11 ),
       .io_out_10( Activation_2_io_out_10 ),
       .io_out_9( Activation_2_io_out_9 ),
       .io_out_8( Activation_2_io_out_8 ),
       .io_out_7( Activation_2_io_out_7 ),
       .io_out_6( Activation_2_io_out_6 ),
       .io_out_5( Activation_2_io_out_5 ),
       .io_out_4( Activation_2_io_out_4 ),
       .io_out_3( Activation_2_io_out_3 ),
       .io_out_2( Activation_2_io_out_2 ),
       .io_out_1( Activation_2_io_out_1 ),
       .io_out_0( Activation_2_io_out_0 )
  );
  MemoryStreamer_1 memoryStreamer(.clk(clk), .reset(reset),
       .io_restart( control_io_memoryRestart ),
       .io_weights_15( memoryStreamer_io_weights_15 ),
       .io_weights_14( memoryStreamer_io_weights_14 ),
       .io_weights_13( memoryStreamer_io_weights_13 ),
       .io_weights_12( memoryStreamer_io_weights_12 ),
       .io_weights_11( memoryStreamer_io_weights_11 ),
       .io_weights_10( memoryStreamer_io_weights_10 ),
       .io_weights_9( memoryStreamer_io_weights_9 ),
       .io_weights_8( memoryStreamer_io_weights_8 ),
       .io_weights_7( memoryStreamer_io_weights_7 ),
       .io_weights_6( memoryStreamer_io_weights_6 ),
       .io_weights_5( memoryStreamer_io_weights_5 ),
       .io_weights_4( memoryStreamer_io_weights_4 ),
       .io_weights_3( memoryStreamer_io_weights_3 ),
       .io_weights_2( memoryStreamer_io_weights_2 ),
       .io_weights_1( memoryStreamer_io_weights_1 ),
       .io_weights_0( memoryStreamer_io_weights_0 ),
       .io_bias( memoryStreamer_io_bias )
  );
endmodule

module MemoryUnit_26(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[7:0] T5;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T6;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (T5)
    0: T0 = 32'h2262841d;
    1: T0 = 32'h499492c2;
    2: T0 = 32'hbc05e444;
    3: T0 = 32'h4ab0632c;
    4: T0 = 32'h373e9e65;
    5: T0 = 32'h91da2164;
    6: T0 = 32'hd87d97cd;
    7: T0 = 32'h5819071;
    8: T0 = 32'h3dbe35e8;
    9: T0 = 32'h862da650;
    10: T0 = 32'ha4c833e1;
    11: T0 = 32'hc876623d;
    12: T0 = 32'h88e53389;
    13: T0 = 32'hed862dbc;
    14: T0 = 32'ha2dd9e90;
    15: T0 = 32'h48be850f;
    16: T0 = 32'h471dd23f;
    17: T0 = 32'h6dc32e9c;
    18: T0 = 32'hf2a96765;
    19: T0 = 32'h9afa800f;
    20: T0 = 32'h26f08dea;
    21: T0 = 32'hfed77652;
    22: T0 = 32'h5bbd6ac9;
    23: T0 = 32'h9237c02c;
    24: T0 = 32'h7613abb1;
    25: T0 = 32'h66e61e79;
    26: T0 = 32'hc80c43d2;
    27: T0 = 32'ha02d488e;
    28: T0 = 32'h7df1c045;
    29: T0 = 32'h7dae7543;
    30: T0 = 32'hd67f365c;
    31: T0 = 32'hb1e10a61;
    32: T0 = 32'h335e6643;
    33: T0 = 32'hdbb6ea39;
    34: T0 = 32'h7c4d93fa;
    35: T0 = 32'h52b968d8;
    36: T0 = 32'hbcbe79f7;
    37: T0 = 32'habda9ebd;
    38: T0 = 32'h5c7aa076;
    39: T0 = 32'h8b37713;
    40: T0 = 32'h2d9f607e;
    41: T0 = 32'hc787cb45;
    42: T0 = 32'h482e9d0e;
    43: T0 = 32'hcd72fdb2;
    44: T0 = 32'h92156dcf;
    45: T0 = 32'hc4469678;
    46: T0 = 32'hb1d385b3;
    47: T0 = 32'h45ad3bda;
    48: T0 = 32'h5e4d9717;
    49: T0 = 32'h3568e2c9;
    50: T0 = 32'h4da2613e;
    51: T0 = 32'h3bc360ad;
    52: T0 = 32'hd5739ffe;
    53: T0 = 32'h4485d21f;
    54: T0 = 32'ha9860881;
    55: T0 = 32'h576e651e;
    56: T0 = 32'h3a6144ef;
    57: T0 = 32'h696e8e6c;
    58: T0 = 32'h23dd5faa;
    59: T0 = 32'h8015d9bd;
    60: T0 = 32'h66626d8e;
    61: T0 = 32'h38390c73;
    62: T0 = 32'ha22c1eee;
    63: T0 = 32'h8857231f;
    64: T0 = 32'hdce00d49;
    65: T0 = 32'h7eb0ada6;
    66: T0 = 32'h9c23ff47;
    67: T0 = 32'h1ab9e730;
    68: T0 = 32'hbf121464;
    69: T0 = 32'hf8526ba5;
    70: T0 = 32'h1dfc754c;
    71: T0 = 32'hd032eb21;
    72: T0 = 32'h1d873ce1;
    73: T0 = 32'h4e16bd4f;
    74: T0 = 32'h75a22221;
    75: T0 = 32'hec6dacde;
    76: T0 = 32'hb2679939;
    77: T0 = 32'h83104e6a;
    78: T0 = 32'h72fe6a16;
    79: T0 = 32'h6921c0eb;
    80: T0 = 32'hd6e669f0;
    81: T0 = 32'h21d99524;
    82: T0 = 32'h7a29ae3;
    83: T0 = 32'hb3c39fb0;
    84: T0 = 32'h9774f24a;
    85: T0 = 32'h404d51fd;
    86: T0 = 32'he1e0352a;
    87: T0 = 32'h276effe3;
    88: T0 = 32'hf2f0e6c1;
    89: T0 = 32'ha8c9b18a;
    90: T0 = 32'h31df806f;
    91: T0 = 32'ha013ac66;
    92: T0 = 32'h6f664d5f;
    93: T0 = 32'h82152ec;
    94: T0 = 32'hb20cf91f;
    95: T0 = 32'he855f75e;
    96: T0 = 32'hc44844ef;
    97: T0 = 32'h70bedbba;
    98: T0 = 32'h2f3b9c80;
    99: T0 = 32'h17b8cad3;
    100: T0 = 32'h89de7ea5;
    101: T0 = 32'he5b02c22;
    102: T0 = 32'hdcfafaf7;
    103: T0 = 32'heaa252ad;
    104: T0 = 32'hbcae515e;
    105: T0 = 32'hdb194355;
    106: T0 = 32'h7b4db299;
    107: T0 = 32'hdadbf330;
    108: T0 = 32'hf07533f8;
    109: T0 = 32'h9240a57e;
    110: T0 = 32'hf54b85e1;
    111: T0 = 32'h5e15da2;
    112: T0 = 32'he6468e8;
    113: T0 = 32'hedb10d26;
    114: T0 = 32'hd2c21bc1;
    115: T0 = 32'ha442df52;
    116: T0 = 32'h76244201;
    117: T0 = 32'hdac5ade2;
    118: T0 = 32'h1154f77a;
    119: T0 = 32'h87449acd;
    120: T0 = 32'h10ddb91f;
    121: T0 = 32'hfecc7197;
    122: T0 = 32'h84fc8055;
    123: T0 = 32'ha04c2262;
    124: T0 = 32'h67659371;
    125: T0 = 32'h7f88e288;
    126: T0 = 32'h9b3c6115;
    127: T0 = 32'hd9fdcce7;
    128: T0 = 32'h251e82f7;
    129: T0 = 32'hdb5162b8;
    130: T0 = 32'hb404c5ec;
    131: T0 = 32'hcc424a8c;
    132: T0 = 32'hb5304cbf;
    133: T0 = 32'h415a0799;
    134: T0 = 32'hc6dbeaa2;
    135: T0 = 32'h11405430;
    136: T0 = 32'h1750b472;
    137: T0 = 32'hca2dcf55;
    138: T0 = 32'hadea7388;
    139: T0 = 32'h8d5e5b93;
    140: T0 = 32'hcfcf75cf;
    141: T0 = 32'hec861d5b;
    142: T0 = 32'h1a1186fa;
    143: T0 = 32'h48be21da;
    144: T0 = 32'hf2983ff8;
    145: T0 = 32'h6fc15556;
    146: T0 = 32'he0a178e1;
    147: T0 = 32'h9babb531;
    148: T0 = 32'h7ab1134a;
    149: T0 = 32'h7ecfd1d6;
    150: T0 = 32'ha9d1556;
    151: T0 = 32'h11be2b8f;
    152: T0 = 32'h7753eecf;
    153: T0 = 32'h6466249e;
    154: T0 = 32'hc98ecc76;
    155: T0 = 32'hac2f2664;
    156: T0 = 32'hbdf0283f;
    157: T0 = 32'h4def9a8c;
    158: T0 = 32'h52294936;
    159: T0 = 32'hf9b3d61f;
    160: T0 = 32'h31da2914;
    161: T0 = 32'heef1bc07;
    162: T0 = 32'h92722674;
    163: T0 = 32'h9ac8b77e;
    164: T0 = 32'h6ed191da;
    165: T0 = 32'h7a11d8ee;
    166: T0 = 32'h2de44103;
    167: T0 = 32'hd2763d3a;
    168: T0 = 32'h16cd87a9;
    169: T0 = 32'h765ea9ca;
    170: T0 = 32'he1334a52;
    171: T0 = 32'hac4d80cd;
    172: T0 = 32'h3663a4a0;
    173: T0 = 32'hffc9a6d3;
    174: T0 = 32'h353448e7;
    175: T0 = 32'hd1b14665;
    176: T0 = 32'hfce60fc5;
    177: T0 = 32'hdad8e0f1;
    178: T0 = 32'h3d55806b;
    179: T0 = 32'h689564b9;
    180: T0 = 32'hbd03fe77;
    181: T0 = 32'ha14a429d;
    182: T0 = 32'hd653b0fd;
    183: T0 = 32'h5d116743;
    184: T0 = 32'h8d8574e6;
    185: T0 = 32'hea97968d;
    186: T0 = 32'h3ca225af;
    187: T0 = 32'h4d564d90;
    188: T0 = 32'h846b4f3f;
    189: T0 = 32'hc111526e;
    190: T0 = 32'h3881bb16;
    191: T0 = 32'h7a1e31da;
    192: T0 = 32'hdaa5d3b6;
    193: T0 = 32'h21be7b0f;
    194: T0 = 32'ha2ab5238;
    195: T0 = 32'h93e0b0fe;
    196: T0 = 32'h12ee279a;
    197: T0 = 32'h5ec7d87a;
    198: T0 = 32'h59cc4833;
    199: T0 = 32'ha6262dae;
    200: T0 = 32'h30eac78a;
    201: T0 = 32'h86c06a2e;
    202: T0 = 32'h531cddf2;
    203: T0 = 32'ha2e990f5;
    204: T0 = 32'h7064a4f2;
    205: T0 = 32'h17e0a1d3;
    206: T0 = 32'hd74f056d;
    207: T0 = 32'ha5c15665;
    208: T0 = 32'h474f174e;
    209: T0 = 32'hf22acbf8;
    210: T0 = 32'h6dbff94e;
    211: T0 = 32'h138948e9;
    212: T0 = 32'h99ce7ea5;
    213: T0 = 32'h65aaae01;
    214: T0 = 32'h8eb3a27e;
    215: T0 = 32'h6c2ae261;
    216: T0 = 32'h9eac516e;
    217: T0 = 32'h89260b15;
    218: T0 = 32'h7b1536a9;
    219: T0 = 32'h96db7798;
    220: T0 = 32'h78d23a7f;
    221: T0 = 32'h60318f28;
    222: T0 = 32'hf248a613;
    223: T0 = 32'h2511f99a;
    224: T0 = 32'h9cf0ec19;
    225: T0 = 32'hd2b78338;
    226: T0 = 32'h4af9ac5e;
    227: T0 = 32'hc4a842c0;
    228: T0 = 32'h6ccb1e65;
    229: T0 = 32'hdcb427a5;
    230: T0 = 32'h1c5be36d;
    231: T0 = 32'heab1d0f1;
    232: T0 = 32'h49f30d0;
    233: T0 = 32'h5f1ff6f3;
    234: T0 = 32'h4e753a09;
    235: T0 = 32'h2cdd4e0e;
    236: T0 = 32'h5331d388;
    237: T0 = 32'h76c26572;
    238: T0 = 32'h9d39b6d1;
    239: T0 = 32'h14b9a563;
    240: T0 = 32'h3fb4dbb2;
    241: T0 = 32'hec996e56;
    242: T0 = 32'hb10713b1;
    243: T0 = 32'haead9d2f;
    244: T0 = 32'h171ca10e;
    245: T0 = 32'hba5a1452;
    246: T0 = 32'h36bc2ef1;
    247: T0 = 32'hd5048c9e;
    248: T0 = 32'hd5a3cb07;
    249: T0 = 32'h34d16531;
    250: T0 = 32'hb42ac65a;
    251: T0 = 32'h49226332;
    252: T0 = 32'h86667051;
    253: T0 = 32'hcb1911c9;
    254: T0 = 32'h70f710fc;
    255: T0 = 32'h73481e5c;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[7:0];
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T6 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_27(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[7:0] T5;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T6;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (T5)
    0: T0 = 32'hbd1c5b90;
    1: T0 = 32'hec796c85;
    2: T0 = 32'h133a53b1;
    3: T0 = 32'h9c58952f;
    4: T0 = 32'he85281ce;
    5: T0 = 32'h52a1525b;
    6: T0 = 32'hada40580;
    7: T0 = 32'hd366fd06;
    8: T0 = 32'h52e9e727;
    9: T0 = 32'h195c1c89;
    10: T0 = 32'h6157c17a;
    11: T0 = 32'hb80de5a4;
    12: T0 = 32'h32574c57;
    13: T0 = 32'hb3d8d2db;
    14: T0 = 32'ha73438be;
    15: T0 = 32'hc5215b5c;
    16: T0 = 32'hc4a29e6a;
    17: T0 = 32'h9fe4517d;
    18: T0 = 32'heec51aab;
    19: T0 = 32'h60a76c81;
    20: T0 = 32'h96abbf31;
    21: T0 = 32'hbc4e668d;
    22: T0 = 32'h591db877;
    23: T0 = 32'h289d6a03;
    24: T0 = 32'h6b037456;
    25: T0 = 32'h66a79c93;
    26: T0 = 32'h941e552d;
    27: T0 = 32'h63a23dd9;
    28: T0 = 32'he5bc5b7f;
    29: T0 = 32'h5c3e40a4;
    30: T0 = 32'h48a3fb29;
    31: T0 = 32'h3e6cb9ca;
    32: T0 = 32'h321f1732;
    33: T0 = 32'hce415a6d;
    34: T0 = 32'h911f40b8;
    35: T0 = 32'hd81b68fb;
    36: T0 = 32'h6451cd9a;
    37: T0 = 32'h7a51d85f;
    38: T0 = 32'h3d2418b7;
    39: T0 = 32'hd9750e1b;
    40: T0 = 32'h43c3466e;
    41: T0 = 32'h74dec9cc;
    42: T0 = 32'h80369def;
    43: T0 = 32'h3c2df1f9;
    44: T0 = 32'h9e73648e;
    45: T0 = 32'h9b1c89b5;
    46: T0 = 32'h4a7201a3;
    47: T0 = 32'hf781179c;
    48: T0 = 32'hf5a26ec8;
    49: T0 = 32'h9909d570;
    50: T0 = 32'hb10c9acb;
    51: T0 = 32'h6d56bc51;
    52: T0 = 32'he5246111;
    53: T0 = 32'h156baeb4;
    54: T0 = 32'he2339176;
    55: T0 = 32'h4109ee85;
    56: T0 = 32'hd130785e;
    57: T0 = 32'h89a9b992;
    58: T0 = 32'hb9c8bc0d;
    59: T0 = 32'h1f96bf63;
    60: T0 = 32'hcdcdfb59;
    61: T0 = 32'h888712a0;
    62: T0 = 32'h6c91d833;
    63: T0 = 32'hea1ef0ce;
    64: T0 = 32'h8031992c;
    65: T0 = 32'hf5ea9542;
    66: T0 = 32'hff06cdf;
    67: T0 = 32'h12cb9723;
    68: T0 = 32'h1e972600;
    69: T0 = 32'hea84e142;
    70: T0 = 32'hfd27e59;
    71: T0 = 32'hbe7e8acd;
    72: T0 = 32'hae84c983;
    73: T0 = 32'h660624ba;
    74: T0 = 32'h551761f6;
    75: T0 = 32'ha4f9226e;
    76: T0 = 32'h3c72103b;
    77: T0 = 32'h7257498e;
    78: T0 = 32'hd16e7b1c;
    79: T0 = 32'h7170f425;
    80: T0 = 32'h78cc1736;
    81: T0 = 32'hfad97d8d;
    82: T0 = 32'ha1345838;
    83: T0 = 32'h1667a1ff;
    84: T0 = 32'h9f05afdc;
    85: T0 = 32'hb15a584a;
    86: T0 = 32'hf63d05b3;
    87: T0 = 32'hf908392b;
    88: T0 = 32'hd5e2c7a6;
    89: T0 = 32'ha9b16b0c;
    90: T0 = 32'hbca3c6fb;
    91: T0 = 32'hdd02f0dd;
    92: T0 = 32'h8c0a24b0;
    93: T0 = 32'hc915abd3;
    94: T0 = 32'h74d30d27;
    95: T0 = 32'hfb1e560d;
    96: T0 = 32'ha8f1e0b8;
    97: T0 = 32'h8dc91b2a;
    98: T0 = 32'hfdc49ac1;
    99: T0 = 32'hec67d346;
    100: T0 = 32'hb6316ac1;
    101: T0 = 32'h90422de4;
    102: T0 = 32'h83cd466;
    103: T0 = 32'h1d9d98ec;
    104: T0 = 32'he3531b54;
    105: T0 = 32'h66e76776;
    106: T0 = 32'hb482a845;
    107: T0 = 32'h6166b266;
    108: T0 = 32'hfaeb378;
    109: T0 = 32'h96fa366;
    110: T0 = 32'h4828e561;
    111: T0 = 32'hda0ec465;
    112: T0 = 32'h709f7eb2;
    113: T0 = 32'h8fbeba5b;
    114: T0 = 32'h7f4b1ab9;
    115: T0 = 32'h5a3d1ed2;
    116: T0 = 32'ha6abfb5a;
    117: T0 = 32'haf5059fd;
    118: T0 = 32'h514cb8b6;
    119: T0 = 32'h18953f8f;
    120: T0 = 32'h88f4646;
    121: T0 = 32'h46c6700e;
    122: T0 = 32'h143acc6f;
    123: T0 = 32'h6976b060;
    124: T0 = 32'ha0641f78;
    125: T0 = 32'h133cd16f;
    126: T0 = 32'h59c765e1;
    127: T0 = 32'h77687ece;
    128: T0 = 32'h770fc685;
    129: T0 = 32'hd4da239;
    130: T0 = 32'ha120c63a;
    131: T0 = 32'hef4748c8;
    132: T0 = 32'hc731fafa;
    133: T0 = 32'h14655e3d;
    134: T0 = 32'heaa5e835;
    135: T0 = 32'h754cd522;
    136: T0 = 32'he2611431;
    137: T0 = 32'h38e1dc23;
    138: T0 = 32'hb9cffd8a;
    139: T0 = 32'h32a59d9b;
    140: T0 = 32'heccbc7ce;
    141: T0 = 32'h993d5c73;
    142: T0 = 32'h4626f5eb;
    143: T0 = 32'heb173bf2;
    144: T0 = 32'hc0a3164f;
    145: T0 = 32'he9b1e2b8;
    146: T0 = 32'h9682e546;
    147: T0 = 32'ha2c040e8;
    148: T0 = 32'h962f44af;
    149: T0 = 32'h9ac6eea1;
    150: T0 = 32'h114c2aef;
    151: T0 = 32'h170cf271;
    152: T0 = 32'h319531b9;
    153: T0 = 32'heecddb55;
    154: T0 = 32'h24aa369a;
    155: T0 = 32'he07c5d9b;
    156: T0 = 32'h226470e7;
    157: T0 = 32'h2788dc68;
    158: T0 = 32'h93ed961a;
    159: T0 = 32'hd9f40998;
    160: T0 = 32'h674f376e;
    161: T0 = 32'hb468295d;
    162: T0 = 32'h8d563b9f;
    163: T0 = 32'hbfc381f3;
    164: T0 = 32'hcd072f30;
    165: T0 = 32'h2b016aa7;
    166: T0 = 32'haca278fe;
    167: T0 = 32'hff7e6a43;
    168: T0 = 32'hcae14146;
    169: T0 = 32'h3951131f;
    170: T0 = 32'h353357b7;
    171: T0 = 32'h7405b4d8;
    172: T0 = 32'h26ca9135;
    173: T0 = 32'h937143ea;
    174: T0 = 32'h66a43701;
    175: T0 = 32'he71178c1;
    176: T0 = 32'he8e13517;
    177: T0 = 32'hda40a1ad;
    178: T0 = 32'h1c54973e;
    179: T0 = 32'h7c49626c;
    180: T0 = 32'hbd137ffb;
    181: T0 = 32'h41125a29;
    182: T0 = 32'hce736182;
    183: T0 = 32'h1150f163;
    184: T0 = 32'h8f949420;
    185: T0 = 32'h4b9fdb0c;
    186: T0 = 32'h29e25283;
    187: T0 = 32'h9d56dcbd;
    188: T0 = 32'h9bcb8d36;
    189: T0 = 32'hed03e65b;
    190: T0 = 32'h28902746;
    191: T0 = 32'h4aaf0bf1;
    192: T0 = 32'hd6942137;
    193: T0 = 32'h972c22a9;
    194: T0 = 32'h194797f8;
    195: T0 = 32'h7d150aec;
    196: T0 = 32'ha13147fe;
    197: T0 = 32'h520509b;
    198: T0 = 32'he922642a;
    199: T0 = 32'hdd61b17e;
    200: T0 = 32'haae897a8;
    201: T0 = 32'hdb854b4c;
    202: T0 = 32'h3792b2fb;
    203: T0 = 32'h51d559a4;
    204: T0 = 32'ha64f44c6;
    205: T0 = 32'h9a79b75b;
    206: T0 = 32'h78ae84d1;
    207: T0 = 32'hab360f68;
    208: T0 = 32'hc4213f48;
    209: T0 = 32'h25c79536;
    210: T0 = 32'he0fd1ac1;
    211: T0 = 32'haaafed72;
    212: T0 = 32'h7eb97341;
    213: T0 = 32'hfe7fe882;
    214: T0 = 32'h728d156e;
    215: T0 = 32'h37fc3a69;
    216: T0 = 32'he7436845;
    217: T0 = 32'h7466e9de;
    218: T0 = 32'h948f8425;
    219: T0 = 32'h25afb4c3;
    220: T0 = 32'hddb8aa3b;
    221: T0 = 32'h5d3fe228;
    222: T0 = 32'h52656917;
    223: T0 = 32'hfa13d4a1;
    224: T0 = 32'h339af257;
    225: T0 = 32'hc0b74af9;
    226: T0 = 32'h5ad9939b;
    227: T0 = 32'hc53c68de;
    228: T0 = 32'h28f79b5;
    229: T0 = 32'h98be1e55;
    230: T0 = 32'h175be8b7;
    231: T0 = 32'hea81169e;
    232: T0 = 32'h81bef71e;
    233: T0 = 32'h955c4b15;
    234: T0 = 32'hc421bcf9;
    235: T0 = 32'h7b883f31;
    236: T0 = 32'h4b38774a;
    237: T0 = 32'h75869563;
    238: T0 = 32'h1d5385e1;
    239: T0 = 32'h92f83bf6;
    240: T0 = 32'h233d24db;
    241: T0 = 32'he8d102b2;
    242: T0 = 32'hc6d0bb42;
    243: T0 = 32'had425b74;
    244: T0 = 32'h7f0c5285;
    245: T0 = 32'hc04eaea5;
    246: T0 = 32'h8493b76e;
    247: T0 = 32'h27f9f270;
    248: T0 = 32'h8674b878;
    249: T0 = 32'hee3da9d4;
    250: T0 = 32'ha9e0a21d;
    251: T0 = 32'h8d5c6fe2;
    252: T0 = 32'h4fef3a89;
    253: T0 = 32'h6cc7863c;
    254: T0 = 32'hba198a17;
    255: T0 = 32'hd89ee1d2;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[7:0];
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T6 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_28(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[7:0] T5;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T6;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (T5)
    0: T0 = 32'h39f073ae;
    1: T0 = 32'h4e472d3c;
    2: T0 = 32'hd3791381;
    3: T0 = 32'hd83a89ce;
    4: T0 = 32'h4cd165b8;
    5: T0 = 32'hbeb1eec2;
    6: T0 = 32'h7f2c6c72;
    7: T0 = 32'h9877dd0c;
    8: T0 = 32'h4e83c930;
    9: T0 = 32'h54567b41;
    10: T0 = 32'hd637969b;
    11: T0 = 32'hff2979d2;
    12: T0 = 32'hb631d071;
    13: T0 = 32'h9f3cf44a;
    14: T0 = 32'h4de70551;
    15: T0 = 32'h7761dcf0;
    16: T0 = 32'h338e923e;
    17: T0 = 32'hf33c794f;
    18: T0 = 32'h1d566c35;
    19: T0 = 32'h7dc5a127;
    20: T0 = 32'hbd66a7fa;
    21: T0 = 32'h108d86a;
    22: T0 = 32'ha4e25191;
    23: T0 = 32'h7500092a;
    24: T0 = 32'h8dbc8fa0;
    25: T0 = 32'h8b097e6a;
    26: T0 = 32'h6d715bd2;
    27: T0 = 32'hcd5780cd;
    28: T0 = 32'h6a4e8078;
    29: T0 = 32'he041ad93;
    30: T0 = 32'hb0802728;
    31: T0 = 32'h61646a5;
    32: T0 = 32'hcc65f938;
    33: T0 = 32'he257bdc6;
    34: T0 = 32'h193a3ae7;
    35: T0 = 32'h9d50baf3;
    36: T0 = 32'he9c62008;
    37: T0 = 32'h40a149c6;
    38: T0 = 32'haeb6157a;
    39: T0 = 32'hd1662aac;
    40: T0 = 32'h92b86302;
    41: T0 = 32'h9958219f;
    42: T0 = 32'heb75e075;
    43: T0 = 32'hba99346e;
    44: T0 = 32'h1ad30839;
    45: T0 = 32'hf3c8120d;
    46: T0 = 32'hae704b55;
    47: T0 = 32'h84a3d48c;
    48: T0 = 32'h8ca2eee3;
    49: T0 = 32'h2586c379;
    50: T0 = 32'ha18b92aa;
    51: T0 = 32'hf3357699;
    52: T0 = 32'h2b87a99;
    53: T0 = 32'hbefd114c;
    54: T0 = 32'h59ac861c;
    55: T0 = 32'h24a6aa97;
    56: T0 = 32'h796b745e;
    57: T0 = 32'h14e0c43b;
    58: T0 = 32'hd20cac69;
    59: T0 = 32'h72ab3370;
    60: T0 = 32'hf0d43f5e;
    61: T0 = 32'h8d3e15ef;
    62: T0 = 32'hc7ebd5e0;
    63: T0 = 32'hb540334e;
    64: T0 = 32'h2b4bf215;
    65: T0 = 32'h132e186a;
    66: T0 = 32'h6dc64c54;
    67: T0 = 32'h71a5e946;
    68: T0 = 32'h99ef45b1;
    69: T0 = 32'h458eac72;
    70: T0 = 32'hc042da60;
    71: T0 = 32'h2fb980bc;
    72: T0 = 32'h280e9b5c;
    73: T0 = 32'h8b2a6bf4;
    74: T0 = 32'h635d1ed0;
    75: T0 = 32'h46da124f;
    76: T0 = 32'h71fcf6c8;
    77: T0 = 32'h30f7ac14;
    78: T0 = 32'hbb0942a1;
    79: T0 = 32'h6168425;
    80: T0 = 32'h5e1d6cd1;
    81: T0 = 32'hf23682b2;
    82: T0 = 32'h5a9f9a4a;
    83: T0 = 32'h13b87ed8;
    84: T0 = 32'ha8ce5ac5;
    85: T0 = 32'he7b005e5;
    86: T0 = 32'hf442936e;
    87: T0 = 32'h4aa132dd;
    88: T0 = 32'h1c3e7658;
    89: T0 = 32'h8b9880d4;
    90: T0 = 32'h427da849;
    91: T0 = 32'h5fd90f67;
    92: T0 = 32'h502d7f8d;
    93: T0 = 32'hb4c0167c;
    94: T0 = 32'hb5c4c8d1;
    95: T0 = 32'h5e9a55e;
    96: T0 = 32'h5e6531b7;
    97: T0 = 32'hcab56ebe;
    98: T0 = 32'h9a0b03c2;
    99: T0 = 32'hc40c59ee;
    100: T0 = 32'h5e0e45ae;
    101: T0 = 32'h9073c293;
    102: T0 = 32'ha77466aa;
    103: T0 = 32'hea01f46e;
    104: T0 = 32'h85dcab29;
    105: T0 = 32'h39997b49;
    106: T0 = 32'h6c6382bb;
    107: T0 = 32'h7d40f9b6;
    108: T0 = 32'hb0f4477;
    109: T0 = 32'he781f74b;
    110: T0 = 32'h3d95a457;
    111: T0 = 32'hd2be09d8;
    112: T0 = 32'ha932eed3;
    113: T0 = 32'hfaeb983b;
    114: T0 = 32'h4cf99c98;
    115: T0 = 32'h938b7cc2;
    116: T0 = 32'h59d3d0b1;
    117: T0 = 32'h69938ef2;
    118: T0 = 32'he91d866;
    119: T0 = 32'haa76969d;
    120: T0 = 32'hd695791f;
    121: T0 = 32'hf07fe963;
    122: T0 = 32'h4b15bc4d;
    123: T0 = 32'hac19bf73;
    124: T0 = 32'h3f12f7c8;
    125: T0 = 32'h5647bc70;
    126: T0 = 32'h5448c4b1;
    127: T0 = 32'h853198b0;
    128: T0 = 32'hb9d86c93;
    129: T0 = 32'he971a4a9;
    130: T0 = 32'h46c282ba;
    131: T0 = 32'hec4268d8;
    132: T0 = 32'h1e35d2fe;
    133: T0 = 32'hd84756bd;
    134: T0 = 32'h1d70023;
    135: T0 = 32'h174c771b;
    136: T0 = 32'h12d5467a;
    137: T0 = 32'heecfc94c;
    138: T0 = 32'h4f0beeb;
    139: T0 = 32'ha140ddb5;
    140: T0 = 32'h4f666dce;
    141: T0 = 32'h7e8f967b;
    142: T0 = 32'h1a2cc5fb;
    143: T0 = 32'hde9e13da;
    144: T0 = 32'hf51e61d7;
    145: T0 = 32'h216fe6b8;
    146: T0 = 32'h63e883ea;
    147: T0 = 32'hb3877acc;
    148: T0 = 32'h42aed6fe;
    149: T0 = 32'haea70edd;
    150: T0 = 32'h6305aaa7;
    151: T0 = 32'h26ca775e;
    152: T0 = 32'hfa61b778;
    153: T0 = 32'hb0604b45;
    154: T0 = 32'h3619a2ca;
    155: T0 = 32'h22b37fb5;
    156: T0 = 32'h65b66cc6;
    157: T0 = 32'h1a779c79;
    158: T0 = 32'hc74e94f1;
    159: T0 = 32'hb3552bde;
    160: T0 = 32'h295bcd91;
    161: T0 = 32'h78a79202;
    162: T0 = 32'h2d3dc874;
    163: T0 = 32'h13bb3630;
    164: T0 = 32'h9c0cd2c3;
    165: T0 = 32'ha97a11fc;
    166: T0 = 32'h5ebb9705;
    167: T0 = 32'h2881379b;
    168: T0 = 32'he52656cc;
    169: T0 = 32'ha0b584ce;
    170: T0 = 32'h7d83a865;
    171: T0 = 32'hd3233365;
    172: T0 = 32'h8d826f8e;
    173: T0 = 32'hc9570ab5;
    174: T0 = 32'h5443d8a4;
    175: T0 = 32'hf53e771e;
    176: T0 = 32'h3bf81526;
    177: T0 = 32'h2cc1ffab;
    178: T0 = 32'ha5b01aba;
    179: T0 = 32'haa4763f3;
    180: T0 = 32'h763137c5;
    181: T0 = 32'h586959ee;
    182: T0 = 32'h63bd0536;
    183: T0 = 32'h974c3a0b;
    184: T0 = 32'he34346c6;
    185: T0 = 32'h7476c39e;
    186: T0 = 32'hb88ed2ef;
    187: T0 = 32'ha524f075;
    188: T0 = 32'hafc312fe;
    189: T0 = 32'hd2fcb6f;
    190: T0 = 32'h4e3c2561;
    191: T0 = 32'hf81e574f;
    192: T0 = 32'hf19ade60;
    193: T0 = 32'he8d95dd4;
    194: T0 = 32'h93e58c0;
    195: T0 = 32'ha747f463;
    196: T0 = 32'h9b0c4105;
    197: T0 = 32'h16a8144;
    198: T0 = 32'hae331f7d;
    199: T0 = 32'h6e680a45;
    200: T0 = 32'hd1606e6f;
    201: T0 = 32'ha93121de;
    202: T0 = 32'h3d630c4d;
    203: T0 = 32'h1b9067d1;
    204: T0 = 32'hce867eef;
    205: T0 = 32'hc3511ba4;
    206: T0 = 32'h6442cac6;
    207: T0 = 32'ha65ef49f;
    208: T0 = 32'h8861e971;
    209: T0 = 32'h2fc246c0;
    210: T0 = 32'hf2e1a046;
    211: T0 = 32'h98ba56a1;
    212: T0 = 32'h68f1c847;
    213: T0 = 32'h7e95a1d7;
    214: T0 = 32'h5b8d174c;
    215: T0 = 32'h907706d4;
    216: T0 = 32'h6e03eecf;
    217: T0 = 32'h566e84f8;
    218: T0 = 32'hc19ea144;
    219: T0 = 32'hb42d6f66;
    220: T0 = 32'hf5f17e8f;
    221: T0 = 32'h3fbe1b2c;
    222: T0 = 32'h8b2fd8d6;
    223: T0 = 32'h9a1f51c;
    224: T0 = 32'h73defec0;
    225: T0 = 32'ha6439435;
    226: T0 = 32'hd3591e8b;
    227: T0 = 32'hd8bffd50;
    228: T0 = 32'h60d14151;
    229: T0 = 32'hfe71aeb3;
    230: T0 = 32'h7f2dd177;
    231: T0 = 32'h9a37c787;
    232: T0 = 32'h4a83697f;
    233: T0 = 32'h54569983;
    234: T0 = 32'hdc179c15;
    235: T0 = 32'hfd299fd3;
    236: T0 = 32'h9411ef5f;
    237: T0 = 32'h9f3e3630;
    238: T0 = 32'h4de6c833;
    239: T0 = 32'h3761d8f0;
    240: T0 = 32'h3fce5ba8;
    241: T0 = 32'hd2496d4c;
    242: T0 = 32'he17972b1;
    243: T0 = 32'h5bbf9d27;
    244: T0 = 32'h4cc1a10a;
    245: T0 = 32'h2539d65b;
    246: T0 = 32'hce1f5c91;
    247: T0 = 32'hb8f30d8e;
    248: T0 = 32'hc607cf2f;
    249: T0 = 32'h6037192b;
    250: T0 = 32'hd913cd5e;
    251: T0 = 32'h1d8e30ae;
    252: T0 = 32'h3d9bc457;
    253: T0 = 32'hd95ff181;
    254: T0 = 32'h5420652e;
    255: T0 = 32'hbc3b5adc;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[7:0];
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T6 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_29(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[7:0] T5;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T6;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (T5)
    0: T0 = 32'h5e1d9e68;
    1: T0 = 32'h2117d17d;
    2: T0 = 32'ha1ad1bbf;
    3: T0 = 32'h173d4c91;
    4: T0 = 32'h2682731;
    5: T0 = 32'h35fa6f1d;
    6: T0 = 32'hca2dba75;
    7: T0 = 32'h40a34a07;
    8: T0 = 32'h732a7456;
    9: T0 = 32'h10201c13;
    10: T0 = 32'hdb0c7d25;
    11: T0 = 32'hd28a3d50;
    12: T0 = 32'hddb95b7f;
    13: T0 = 32'h8df644a6;
    14: T0 = 32'he75bfb09;
    15: T0 = 32'h254679ca;
    16: T0 = 32'h362e851;
    17: T0 = 32'h70684694;
    18: T0 = 32'h2d3e8dc6;
    19: T0 = 32'h37457f8c;
    20: T0 = 32'hc946c0ce;
    21: T0 = 32'h412886d3;
    22: T0 = 32'haea21708;
    23: T0 = 32'hf86a97d4;
    24: T0 = 32'hcb64af39;
    25: T0 = 32'ha93129e1;
    26: T0 = 32'h3ba3ac5c;
    27: T0 = 32'h17944f83;
    28: T0 = 32'hae8a6e87;
    29: T0 = 32'hc251ba18;
    30: T0 = 32'h60c0d8fe;
    31: T0 = 32'h261fbc1c;
    32: T0 = 32'hc0e13e4a;
    33: T0 = 32'hc6b7c17d;
    34: T0 = 32'h4afd1abf;
    35: T0 = 32'h47fc4c91;
    36: T0 = 32'h488f7f31;
    37: T0 = 32'h6eb3679d;
    38: T0 = 32'h155db875;
    39: T0 = 32'haab56e87;
    40: T0 = 32'h4966476;
    41: T0 = 32'hda5e94b7;
    42: T0 = 32'h4631742c;
    43: T0 = 32'h7de09dd8;
    44: T0 = 32'hb39597e;
    45: T0 = 32'h76cb50a6;
    46: T0 = 32'h9d74ff03;
    47: T0 = 32'h76ea79ca;
    48: T0 = 32'h3b9a1317;
    49: T0 = 32'hdb246ae8;
    50: T0 = 32'h7d5d4554;
    51: T0 = 32'h5bb169ee;
    52: T0 = 32'h9d2747a5;
    53: T0 = 32'ha10a9842;
    54: T0 = 32'hd85b08a7;
    55: T0 = 32'h3831201b;
    56: T0 = 32'h2f8edd6e;
    57: T0 = 32'hcfa74b54;
    58: T0 = 32'h3d3b3eda;
    59: T0 = 32'hcd72f7b9;
    60: T0 = 32'hb14034ee;
    61: T0 = 32'hc053ad1d;
    62: T0 = 32'hf0c906e6;
    63: T0 = 32'h752e0db9;
    64: T0 = 32'h5ed496a4;
    65: T0 = 32'hde01db49;
    66: T0 = 32'hb05dc83d;
    67: T0 = 32'h6c3d6491;
    68: T0 = 32'ha401bf31;
    69: T0 = 32'hf1305d5c;
    70: T0 = 32'hb67d9a95;
    71: T0 = 32'hd8150c8f;
    72: T0 = 32'h859f56d6;
    73: T0 = 32'h569f8636;
    74: T0 = 32'hace27da0;
    75: T0 = 32'h5d442239;
    76: T0 = 32'h9e1b9fbe;
    77: T0 = 32'he5824da7;
    78: T0 = 32'h28b03768;
    79: T0 = 32'h5eae3f8f;
    80: T0 = 32'h12a37ec8;
    81: T0 = 32'hf26a9d26;
    82: T0 = 32'h6dbe1ad3;
    83: T0 = 32'h13c1bd72;
    84: T0 = 32'h89ce3140;
    85: T0 = 32'h67a8a8a6;
    86: T0 = 32'hebd2d572;
    87: T0 = 32'h6c72bbc1;
    88: T0 = 32'hbc0c4997;
    89: T0 = 32'hcb313187;
    90: T0 = 32'h7b558c05;
    91: T0 = 32'h96db9a63;
    92: T0 = 32'h78d2c331;
    93: T0 = 32'hd031e2c2;
    94: T0 = 32'hf34a6d13;
    95: T0 = 32'h2471cce4;
    96: T0 = 32'hd8f08579;
    97: T0 = 32'h836e46d6;
    98: T0 = 32'h66d5e046;
    99: T0 = 32'he04f4609;
    100: T0 = 32'h41ed8c07;
    101: T0 = 32'h4fa72305;
    102: T0 = 32'h631b3fcd;
    103: T0 = 32'h3a9d42d1;
    104: T0 = 32'h4e4e3cdf;
    105: T0 = 32'heb6e86f1;
    106: T0 = 32'h877d2304;
    107: T0 = 32'hf9c6fee;
    108: T0 = 32'h6db97aaf;
    109: T0 = 32'h7a7f18ac;
    110: T0 = 32'h9d80da9e;
    111: T0 = 32'h1a3aa19b;
    112: T0 = 32'h3b9904e7;
    113: T0 = 32'h116f62f8;
    114: T0 = 32'h2dbca1ce;
    115: T0 = 32'ha7e74aad;
    116: T0 = 32'h43aedea7;
    117: T0 = 32'h2caf6787;
    118: T0 = 32'he20baefc;
    119: T0 = 32'h2ecbe661;
    120: T0 = 32'hf1626472;
    121: T0 = 32'ha1a0d315;
    122: T0 = 32'h5b4923ae;
    123: T0 = 32'h129a6dba;
    124: T0 = 32'h75925e6f;
    125: T0 = 32'h40775a2c;
    126: T0 = 32'hf64bb058;
    127: T0 = 32'ha75f299a;
    128: T0 = 32'h9798017;
    129: T0 = 32'h337766c9;
    130: T0 = 32'h6cb8c56e;
    131: T0 = 32'h13c0428f;
    132: T0 = 32'h1beeceb6;
    133: T0 = 32'h458e5119;
    134: T0 = 32'hca932e8d;
    135: T0 = 32'h262ac43f;
    136: T0 = 32'hf060d4a8;
    137: T0 = 32'ha121c671;
    138: T0 = 32'h5b4d33fa;
    139: T0 = 32'h8a9b6b9c;
    140: T0 = 32'h69b26486;
    141: T0 = 32'h60759d7d;
    142: T0 = 32'hd64b96f8;
    143: T0 = 32'ha457231c;
    144: T0 = 32'h958f8b1;
    145: T0 = 32'h6cd1de72;
    146: T0 = 32'h92a2cc78;
    147: T0 = 32'h8a48fd82;
    148: T0 = 32'h7ed8c090;
    149: T0 = 32'hdaf5a552;
    150: T0 = 32'h25e4da15;
    151: T0 = 32'hb76e949e;
    152: T0 = 32'h93f1df1f;
    153: T0 = 32'h365fe460;
    154: T0 = 32'hc1d4ad5c;
    155: T0 = 32'ha84d1367;
    156: T0 = 32'h2e65f680;
    157: T0 = 32'h7f8f3931;
    158: T0 = 32'h67dc0b8;
    159: T0 = 32'hc8f19e34;
    160: T0 = 32'ha15e936e;
    161: T0 = 32'h85376d4d;
    162: T0 = 32'he2d9493d;
    163: T0 = 32'hc57c8127;
    164: T0 = 32'h62a9253a;
    165: T0 = 32'hdebfd81a;
    166: T0 = 32'h525d7c91;
    167: T0 = 32'h2a81cc0e;
    168: T0 = 32'h447681a3;
    169: T0 = 32'h367d3f3b;
    170: T0 = 32'h6755796;
    171: T0 = 32'h63caf09a;
    172: T0 = 32'h6b9d8072;
    173: T0 = 32'h76c6a9c2;
    174: T0 = 32'h9d3d276e;
    175: T0 = 32'h96fa4aa1;
    176: T0 = 32'h2b1c4e41;
    177: T0 = 32'h936c802d;
    178: T0 = 32'h6d5c5e2a;
    179: T0 = 32'h72bde970;
    180: T0 = 32'h910351eb;
    181: T0 = 32'ha93adebd;
    182: T0 = 32'h565b556e;
    183: T0 = 32'h7891f73b;
    184: T0 = 32'hcf0e1079;
    185: T0 = 32'hcf27ebc5;
    186: T0 = 32'h342b9e8d;
    187: T0 = 32'h4fd2fdc1;
    188: T0 = 32'ha19aa6ea;
    189: T0 = 32'hc077a673;
    190: T0 = 32'h59c3cca3;
    191: T0 = 32'h3f2ec8f2;
    192: T0 = 32'h7ad92dee;
    193: T0 = 32'h916ee5a5;
    194: T0 = 32'h4bdab3a3;
    195: T0 = 32'h794512b8;
    196: T0 = 32'h802fbf4a;
    197: T0 = 32'h2f04539d;
    198: T0 = 32'h71023cfa;
    199: T0 = 32'haeda6b47;
    200: T0 = 32'h8cc24a6;
    201: T0 = 32'hb996948f;
    202: T0 = 32'h163be1aa;
    203: T0 = 32'h47f52da0;
    204: T0 = 32'h422a093f;
    205: T0 = 32'h103143cf;
    206: T0 = 32'h51aeb95e;
    207: T0 = 32'h37483bde;
    208: T0 = 32'hfc456d90;
    209: T0 = 32'h924eb403;
    210: T0 = 32'h61dd9aa2;
    211: T0 = 32'h753d3f30;
    212: T0 = 32'h60c5f04a;
    213: T0 = 32'h7bb51fc;
    214: T0 = 32'hee0b1526;
    215: T0 = 32'hc8d139b3;
    216: T0 = 32'h4e2a2644;
    217: T0 = 32'hd9f0a08e;
    218: T0 = 32'h5bb5a06d;
    219: T0 = 32'h5fb2ac64;
    220: T0 = 32'hc999cdc9;
    221: T0 = 32'h903653ff;
    222: T0 = 32'h6d82e9e5;
    223: T0 = 32'ha60a675e;
    224: T0 = 32'h13b14c51;
    225: T0 = 32'hee3ab03d;
    226: T0 = 32'h1b8ac43a;
    227: T0 = 32'hfc446e10;
    228: T0 = 32'he7d6d07b;
    229: T0 = 32'hc205963d;
    230: T0 = 32'hade2910d;
    231: T0 = 32'hd7767733;
    232: T0 = 32'h10fc34f1;
    233: T0 = 32'h5bde88c2;
    234: T0 = 32'h64763d28;
    235: T0 = 32'h3a45cd99;
    236: T0 = 32'h1267cf8f;
    237: T0 = 32'hb2884e73;
    238: T0 = 32'ha93cfa9a;
    239: T0 = 32'h47e123ba;
    240: T0 = 32'hd4271136;
    241: T0 = 32'h13ae6e88;
    242: T0 = 32'h6dc42330;
    243: T0 = 32'h71b192ae;
    244: T0 = 32'h99ef8ece;
    245: T0 = 32'h78e59da;
    246: T0 = 32'hd1c26483;
    247: T0 = 32'h67b23d7e;
    248: T0 = 32'h280e9fa8;
    249: T0 = 32'h8b2f6e4c;
    250: T0 = 32'h63fd42db;
    251: T0 = 32'h6db51bc;
    252: T0 = 32'h61b964c2;
    253: T0 = 32'h3077b55b;
    254: T0 = 32'hbb0805ec;
    255: T0 = 32'h677073d;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[7:0];
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T6 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_30(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[7:0] T5;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T6;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (T5)
    0: T0 = 32'h700f8d2e;
    1: T0 = 32'hdeb7edc5;
    2: T0 = 32'h5e7960af;
    3: T0 = 32'h49816ab;
    4: T0 = 32'hfccfbc4e;
    5: T0 = 32'hccb44019;
    6: T0 = 32'hc530d91;
    7: T0 = 32'h8ab76903;
    8: T0 = 32'h49f66a7;
    9: T0 = 32'h5f1e9489;
    10: T0 = 32'h4e716166;
    11: T0 = 32'hfd49e5ac;
    12: T0 = 32'h5335083e;
    13: T0 = 32'h76ce58ef;
    14: T0 = 32'hbd117a5c;
    15: T0 = 32'h54f13b5f;
    16: T0 = 32'h3f9c1337;
    17: T0 = 32'h6cf16e8b;
    18: T0 = 32'hd2f05178;
    19: T0 = 32'h98c061fa;
    20: T0 = 32'hfe514ea5;
    21: T0 = 32'h5a959942;
    22: T0 = 32'h2dc502b7;
    23: T0 = 32'h937e3a5e;
    24: T0 = 32'h32d5532e;
    25: T0 = 32'h785e4354;
    26: T0 = 32'hc1d4bed9;
    27: T0 = 32'ha44d73b5;
    28: T0 = 32'h367136c8;
    29: T0 = 32'h3fa9af3d;
    30: T0 = 32'h8a3c04e7;
    31: T0 = 32'hc9b15f1f;
    32: T0 = 32'hf59ecb71;
    33: T0 = 32'h9a5156e4;
    34: T0 = 32'hf44484c0;
    35: T0 = 32'h6d767f3c;
    36: T0 = 32'h7585c08e;
    37: T0 = 32'h817e8653;
    38: T0 = 32'hf69f2749;
    39: T0 = 32'h1d19d6d4;
    40: T0 = 32'hc531ab3d;
    41: T0 = 32'h28a929f1;
    42: T0 = 32'h9dca8d5e;
    43: T0 = 32'hf164fef;
    44: T0 = 32'hcd896ec5;
    45: T0 = 32'hed861a11;
    46: T0 = 32'he91c896;
    47: T0 = 32'hda9e809c;
    48: T0 = 32'ha3993641;
    49: T0 = 32'h9604a1bc;
    50: T0 = 32'hf90ded46;
    51: T0 = 32'h6c1cec50;
    52: T0 = 32'he14355ef;
    53: T0 = 32'h15b0aeb5;
    54: T0 = 32'hfc62416a;
    55: T0 = 32'h48d5f371;
    56: T0 = 32'h12b31b1;
    57: T0 = 32'h19fbfbc4;
    58: T0 = 32'hab641f96;
    59: T0 = 32'h5f80cd9b;
    60: T0 = 32'hd89d8c77;
    61: T0 = 32'ha7ba6e52;
    62: T0 = 32'h6cb0ae1e;
    63: T0 = 32'heae89b1;
    64: T0 = 32'hc6a1ee11;
    65: T0 = 32'he2b3903d;
    66: T0 = 32'h22b8cd3e;
    67: T0 = 32'h86ba6f18;
    68: T0 = 32'h5eccd17b;
    69: T0 = 32'hdafaae3d;
    70: T0 = 32'h16fdf800;
    71: T0 = 32'haa22d533;
    72: T0 = 32'h97be1491;
    73: T0 = 32'h9019f8e2;
    74: T0 = 32'hc7737d00;
    75: T0 = 32'hab598e8b;
    76: T0 = 32'h5d36cfcc;
    77: T0 = 32'h6dc67c73;
    78: T0 = 32'hb453f79a;
    79: T0 = 32'h5f9a8f2;
    80: T0 = 32'h2b5aecd1;
    81: T0 = 32'ha45992b3;
    82: T0 = 32'h8282a3ca;
    83: T0 = 32'ha44e5ed8;
    84: T0 = 32'h42d0dae5;
    85: T0 = 32'h5ef50df4;
    86: T0 = 32'h21a4836e;
    87: T0 = 32'hf7ecb7f4;
    88: T0 = 32'hd271725c;
    89: T0 = 32'h30f080d6;
    90: T0 = 32'ha2c4a02d;
    91: T0 = 32'h32a84774;
    92: T0 = 32'h4e1d7f8f;
    93: T0 = 32'h3ba9127c;
    94: T0 = 32'hf3ed9b1;
    95: T0 = 32'h8ad1295e;
    96: T0 = 32'ha1a39647;
    97: T0 = 32'heceb933b;
    98: T0 = 32'h9b3adc3e;
    99: T0 = 32'h9c486850;
    100: T0 = 32'heed277b5;
    101: T0 = 32'h52b5ff64;
    102: T0 = 32'hada4d877;
    103: T0 = 32'hd66e6a23;
    104: T0 = 32'h12fd5456;
    105: T0 = 32'h795dca17;
    106: T0 = 32'he3777ea9;
    107: T0 = 32'hb80d94d9;
    108: T0 = 32'hba6393bc;
    109: T0 = 32'hb3994d76;
    110: T0 = 32'haf242761;
    111: T0 = 32'h81c1bba3;
    112: T0 = 32'hd4a68367;
    113: T0 = 32'hfa9966d8;
    114: T0 = 32'hb557e56e;
    115: T0 = 32'hafa31aad;
    116: T0 = 32'h97158eaf;
    117: T0 = 32'ha15a421b;
    118: T0 = 32'hd6bf2add;
    119: T0 = 32'hfd084654;
    120: T0 = 32'hd5e0e06e;
    121: T0 = 32'ha8919eb9;
    122: T0 = 32'hbca32396;
    123: T0 = 32'h5d124db8;
    124: T0 = 32'h8d0f7cc7;
    125: T0 = 32'hc9171c8c;
    126: T0 = 32'h60d39ada;
    127: T0 = 32'hfe1e3998;
    128: T0 = 32'he8f09f41;
    129: T0 = 32'hdac0e495;
    130: T0 = 32'h1c556d66;
    131: T0 = 32'h7cbdf501;
    132: T0 = 32'hfd53917a;
    133: T0 = 32'hc10ae21b;
    134: T0 = 32'h9ef31501;
    135: T0 = 32'h1910c571;
    136: T0 = 32'hf1da8b9;
    137: T0 = 32'heb9fbdea;
    138: T0 = 32'ha9e21d16;
    139: T0 = 32'hdd540d8b;
    140: T0 = 32'h8b43ec87;
    141: T0 = 32'he4871811;
    142: T0 = 32'h3890da9e;
    143: T0 = 32'h4abeb39b;
    144: T0 = 32'hd0b46099;
    145: T0 = 32'h9317b32a;
    146: T0 = 32'he4cdaf4c;
    147: T0 = 32'hc03e868c;
    148: T0 = 32'h20a9ba61;
    149: T0 = 32'h9ff335a4;
    150: T0 = 32'h521de34c;
    151: T0 = 32'h8995f1a0;
    152: T0 = 32'h453fb090;
    153: T0 = 32'hc4ecf423;
    154: T0 = 32'hce2c7200;
    155: T0 = 32'h7fe20266;
    156: T0 = 32'h7d9d9309;
    157: T0 = 32'h6d8667ce;
    158: T0 = 32'h1dd3f750;
    159: T0 = 32'h9eeaa463;
    160: T0 = 32'h231a1397;
    161: T0 = 32'h60bff281;
    162: T0 = 32'habbbc438;
    163: T0 = 32'hb71f38f8;
    164: T0 = 32'h28edefe;
    165: T0 = 32'hbab0585f;
    166: T0 = 32'h77ac05b1;
    167: T0 = 32'heeee351e;
    168: T0 = 32'hf0e4c60c;
    169: T0 = 32'h34c0c8cc;
    170: T0 = 32'h56119f7b;
    171: T0 = 32'h63a9d1b5;
    172: T0 = 32'h66586;
    173: T0 = 32'h13589b33;
    174: T0 = 32'hd56f19ec;
    175: T0 = 32'hb741271c;
    176: T0 = 32'h2166e4b7;
    177: T0 = 32'hc01382d9;
    178: T0 = 32'hdea2862e;
    179: T0 = 32'hc5444a89;
    180: T0 = 32'h63ecfaf5;
    181: T0 = 32'hc0e737ad;
    182: T0 = 32'h84f2aafc;
    183: T0 = 32'h412050d5;
    184: T0 = 32'h11783454;
    185: T0 = 32'h9ff95631;
    186: T0 = 32'h6bc433a8;
    187: T0 = 32'h2ac87f36;
    188: T0 = 32'h53ad5f8d;
    189: T0 = 32'he68055ef;
    190: T0 = 32'hae10b7f1;
    191: T0 = 32'h88f72b4e;
    192: T0 = 32'h85352998;
    193: T0 = 32'h50eb12e;
    194: T0 = 32'ha389bb73;
    195: T0 = 32'hb3b6e2f0;
    196: T0 = 32'h2f8326b;
    197: T0 = 32'h3eff79ac;
    198: T0 = 32'h59ac450c;
    199: T0 = 32'h24ef7163;
    200: T0 = 32'h792b34c0;
    201: T0 = 32'h4e0ba8e;
    202: T0 = 32'hf60f72a3;
    203: T0 = 32'h73a3c4e5;
    204: T0 = 32'hf0bc8b38;
    205: T0 = 32'hd3c67f3;
    206: T0 = 32'hc7efab41;
    207: T0 = 32'h2544c563;
    208: T0 = 32'h234b148e;
    209: T0 = 32'h3192296b;
    210: T0 = 32'ha8a93abd;
    211: T0 = 32'h83b0a0fa;
    212: T0 = 32'ha3fe3ff0;
    213: T0 = 32'h71de7b6c;
    214: T0 = 32'hdabdd8b6;
    215: T0 = 32'h4522fa8b;
    216: T0 = 32'h753a14c2;
    217: T0 = 32'h8720521e;
    218: T0 = 32'hfbcc53a1;
    219: T0 = 32'hd6ebb018;
    220: T0 = 32'h91d59338;
    221: T0 = 32'h84f665ef;
    222: T0 = 32'he25b3741;
    223: T0 = 32'h25e55fe3;
    224: T0 = 32'h242eeeb;
    225: T0 = 32'h7d1211b6;
    226: T0 = 32'hb02b9d43;
    227: T0 = 32'h9af24dd1;
    228: T0 = 32'ha7704025;
    229: T0 = 32'h50c8aca2;
    230: T0 = 32'h49ecf77e;
    231: T0 = 32'h4506e2d5;
    232: T0 = 32'h3123795e;
    233: T0 = 32'hea161d3;
    234: T0 = 32'he1cc341d;
    235: T0 = 32'ha0213e52;
    236: T0 = 32'hb045fbd9;
    237: T0 = 32'h8db82628;
    238: T0 = 32'he67fc013;
    239: T0 = 32'h6987dca0;
    240: T0 = 32'hc567c2cf;
    241: T0 = 32'h8dd96179;
    242: T0 = 32'he644c18f;
    243: T0 = 32'hece7d8cd;
    244: T0 = 32'hb633ef31;
    245: T0 = 32'h904aa617;
    246: T0 = 32'h402daaf4;
    247: T0 = 32'h1f19c64c;
    248: T0 = 32'hcb51f077;
    249: T0 = 32'h6687db35;
    250: T0 = 32'hb48a1f9a;
    251: T0 = 32'h61466d9a;
    252: T0 = 32'h56cc27f;
    253: T0 = 32'h90e7c08;
    254: T0 = 32'h58a5b719;
    255: T0 = 32'h7a1e3992;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[7:0];
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T6 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_31(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[7:0] T5;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T6;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (T5)
    0: T0 = 32'hc4457f41;
    1: T0 = 32'h960ca4a4;
    2: T0 = 32'h195fcfc2;
    3: T0 = 32'h6c1c7d50;
    4: T0 = 32'he14351cb;
    5: T0 = 32'h15b1cebd;
    6: T0 = 32'hae6b1528;
    7: T0 = 32'hd981f753;
    8: T0 = 32'h129a83c;
    9: T0 = 32'h11bba9c4;
    10: T0 = 32'ha8e28c0e;
    11: T0 = 32'h5d80fdf3;
    12: T0 = 32'h92dfcdef;
    13: T0 = 32'ha3a85651;
    14: T0 = 32'h6cb2c89e;
    15: T0 = 32'h4e8b81da;
    16: T0 = 32'hc6217698;
    17: T0 = 32'h73a0b92b;
    18: T0 = 32'hb92f1fb9;
    19: T0 = 32'h16b9ad56;
    20: T0 = 32'ha9fef172;
    21: T0 = 32'h61faacfa;
    22: T0 = 32'hdcfaf522;
    23: T0 = 32'h40a2bdaa;
    24: T0 = 32'hbd0e9b99;
    25: T0 = 32'h9702f966;
    26: T0 = 32'h7b0790f5;
    27: T0 = 32'hdc7bba67;
    28: T0 = 32'hb0d1a210;
    29: T0 = 32'h8450b653;
    30: T0 = 32'he353652f;
    31: T0 = 32'h256146e1;
    32: T0 = 32'h5e64edb1;
    33: T0 = 32'hce901682;
    34: T0 = 32'h9342a440;
    35: T0 = 32'hd89876bd;
    36: T0 = 32'hbe13d8c7;
    37: T0 = 32'hb01111c0;
    38: T0 = 32'h9df48764;
    39: T0 = 32'h991410d4;
    40: T0 = 32'h1e9d7edc;
    41: T0 = 32'h4e5f84f4;
    42: T0 = 32'h84f6216c;
    43: T0 = 32'h6c656665;
    44: T0 = 32'h12657f8a;
    45: T0 = 32'hbf889bbd;
    46: T0 = 32'hab4d8d0;
    47: T0 = 32'h49a8371e;
    48: T0 = 32'hf6aed238;
    49: T0 = 32'hdab73f4e;
    50: T0 = 32'h5a736554;
    51: T0 = 32'h84bc810f;
    52: T0 = 32'h78cf8130;
    53: T0 = 32'hcbbffd62;
    54: T0 = 32'h1c5aca81;
    55: T0 = 32'haab388bc;
    56: T0 = 32'h49e9b99;
    57: T0 = 32'h575e7671;
    58: T0 = 32'h47755bd2;
    59: T0 = 32'h14d8020f;
    60: T0 = 32'h1b31b290;
    61: T0 = 32'h76c6ad96;
    62: T0 = 32'hb915074c;
    63: T0 = 32'h16b9ce25;
    64: T0 = 32'hbe9cfbba;
    65: T0 = 32'h3e114ed7;
    66: T0 = 32'he4351381;
    67: T0 = 32'h652e9ea7;
    68: T0 = 32'h7510ba0e;
    69: T0 = 32'hc16e1552;
    70: T0 = 32'hc61dae90;
    71: T0 = 32'h11080e8c;
    72: T0 = 32'hc573ef06;
    73: T0 = 32'ha8bb043f;
    74: T0 = 32'h89c0e17f;
    75: T0 = 32'h5d162362;
    76: T0 = 32'h8d8b7251;
    77: T0 = 32'heca7918e;
    78: T0 = 32'hab151f4;
    79: T0 = 32'hda9e7cdc;
    80: T0 = 32'he3983b48;
    81: T0 = 32'hf8f17546;
    82: T0 = 32'h8e367ad1;
    83: T0 = 32'h5c4b575;
    84: T0 = 32'hfc0e0508;
    85: T0 = 32'hc042e9c2;
    86: T0 = 32'ha6531572;
    87: T0 = 32'hfa402ac8;
    88: T0 = 32'h95dccbcf;
    89: T0 = 32'hfb1d25de;
    90: T0 = 32'h6df0c875;
    91: T0 = 32'had5ca045;
    92: T0 = 32'hf0f2830;
    93: T0 = 32'he6c1828c;
    94: T0 = 32'h30116a07;
    95: T0 = 32'hd8bed44d;
    96: T0 = 32'hacf0a1be;
    97: T0 = 32'h802e33c2;
    98: T0 = 32'h53cbe474;
    99: T0 = 32'hf41c96ac;
    100: T0 = 32'h608fae5e;
    101: T0 = 32'hae35514a;
    102: T0 = 32'h25402f89;
    103: T0 = 32'headf18e4;
    104: T0 = 32'h8cd8780;
    105: T0 = 32'h5dda36ba;
    106: T0 = 32'hc63563e0;
    107: T0 = 32'h77b1422c;
    108: T0 = 32'h22191890;
    109: T0 = 32'hb398598f;
    110: T0 = 32'h8da61acc;
    111: T0 = 32'h9760660f;
    112: T0 = 32'h3d27912e;
    113: T0 = 32'h6c914bda;
    114: T0 = 32'hb0213205;
    115: T0 = 32'h8b7a80af;
    116: T0 = 32'h7e70ad34;
    117: T0 = 32'h50ff3142;
    118: T0 = 32'h8ebd7ad9;
    119: T0 = 32'h852488cc;
    120: T0 = 32'hf733db87;
    121: T0 = 32'h3679363b;
    122: T0 = 32'ha9c45714;
    123: T0 = 32'ha86e221a;
    124: T0 = 32'h9dc11231;
    125: T0 = 32'hedce598c;
    126: T0 = 32'ha6513740;
    127: T0 = 32'hc8affc2d;
    128: T0 = 32'h43da5249;
    129: T0 = 32'h83b6edbc;
    130: T0 = 32'h6cf059c2;
    131: T0 = 32'h83a0e952;
    132: T0 = 32'h1f2e45a5;
    133: T0 = 32'h898eaea3;
    134: T0 = 32'h41dad17e;
    135: T0 = 32'h2e8ae251;
    136: T0 = 32'h85de7979;
    137: T0 = 32'heb2feb55;
    138: T0 = 32'h7f09969f;
    139: T0 = 32'h835effdb;
    140: T0 = 32'h6da6e6e9;
    141: T0 = 32'h6447ae20;
    142: T0 = 32'h904d8c93;
    143: T0 = 32'h58fec8b0;
    144: T0 = 32'h3b5c68f8;
    145: T0 = 32'h53ce0ba2;
    146: T0 = 32'h6d3d97c3;
    147: T0 = 32'h1bb99f54;
    148: T0 = 32'hb9f68040;
    149: T0 = 32'h65b825e2;
    150: T0 = 32'hcebbf76a;
    151: T0 = 32'h70b2d1f4;
    152: T0 = 32'hff0eb990;
    153: T0 = 32'hc9373582;
    154: T0 = 32'h7b0f8051;
    155: T0 = 32'hdc9b0e66;
    156: T0 = 32'hf9c14351;
    157: T0 = 32'hc0707648;
    158: T0 = 32'he642e855;
    159: T0 = 32'h2d27e862;
    160: T0 = 32'hdaf00107;
    161: T0 = 32'h6851a12d;
    162: T0 = 32'h92a65736;
    163: T0 = 32'ha742097e;
    164: T0 = 32'h6ee836fa;
    165: T0 = 32'h56a55aad;
    166: T0 = 32'hada46182;
    167: T0 = 32'hc76e7122;
    168: T0 = 32'h70709421;
    169: T0 = 32'h3058db8f;
    170: T0 = 32'he1c4d3aa;
    171: T0 = 32'hb009d999;
    172: T0 = 32'h7a658576;
    173: T0 = 32'h3f88e753;
    174: T0 = 32'ha63c2743;
    175: T0 = 32'hc8d103e3;
    176: T0 = 32'ha552c0b7;
    177: T0 = 32'h7d902e8b;
    178: T0 = 32'hb92b6534;
    179: T0 = 32'h1b7283ae;
    180: T0 = 32'hb770acfa;
    181: T0 = 32'h52c8536a;
    182: T0 = 32'h9ec6a81;
    183: T0 = 32'h556a913c;
    184: T0 = 32'hb1ab9381;
    185: T0 = 32'h2a97629;
    186: T0 = 32'he1ce53d2;
    187: T0 = 32'ha06b400e;
    188: T0 = 32'h9c65c480;
    189: T0 = 32'h8db8fdd3;
    190: T0 = 32'he6ffb7cc;
    191: T0 = 32'h69c70a25;
    192: T0 = 32'h44662117;
    193: T0 = 32'hdbbee2a8;
    194: T0 = 32'h6c778572;
    195: T0 = 32'h32a16bec;
    196: T0 = 32'h9daf46a5;
    197: T0 = 32'ha90aee3d;
    198: T0 = 32'h14daa2a6;
    199: T0 = 32'h2e90f47a;
    200: T0 = 32'h8c8cb538;
    201: T0 = 32'heb1fcb5d;
    202: T0 = 32'h7d39b689;
    203: T0 = 32'hcd5b79b5;
    204: T0 = 32'h733276cf;
    205: T0 = 32'h6853a77b;
    206: T0 = 32'h910984f1;
    207: T0 = 32'h50fc0510;
    208: T0 = 32'h9efc7119;
    209: T0 = 32'h841f2ca6;
    210: T0 = 32'h135a6740;
    211: T0 = 32'hec5cb52e;
    212: T0 = 32'he10181ce;
    213: T0 = 32'he3180d2;
    214: T0 = 32'had41474a;
    215: T0 = 32'hdb5ebd7c;
    216: T0 = 32'h8e9aba9;
    217: T0 = 32'h1dd83dc8;
    218: T0 = 32'ha67283d3;
    219: T0 = 32'h7cc46bce;
    220: T0 = 32'h20e64d1;
    221: T0 = 32'hb388b288;
    222: T0 = 32'h2da4cade;
    223: T0 = 32'h9740cc50;
    224: T0 = 32'h8423c891;
    225: T0 = 32'h952cb625;
    226: T0 = 32'h6dc1cc30;
    227: T0 = 32'h61d73f70;
    228: T0 = 32'h92afc0ca;
    229: T0 = 32'hae0f987d;
    230: T0 = 32'h41421505;
    231: T0 = 32'h1f9d159a;
    232: T0 = 32'h4ac627bd;
    233: T0 = 32'hceeac8cc;
    234: T0 = 32'h16b8a94e;
    235: T0 = 32'h41f48b6d;
    236: T0 = 32'h606ced86;
    237: T0 = 32'h1a343a31;
    238: T0 = 32'hd9acc8be;
    239: T0 = 32'h3f4c0714;
    240: T0 = 32'h6c0d7fe0;
    241: T0 = 32'h3b38bd64;
    242: T0 = 32'h3c261ac3;
    243: T0 = 32'h2670b472;
    244: T0 = 32'hb524710a;
    245: T0 = 32'h14ac9d5;
    246: T0 = 32'hc8fa1576;
    247: T0 = 32'h15026fc1;
    248: T0 = 32'hbd386e2f;
    249: T0 = 32'haba9098e;
    250: T0 = 32'hb9caa465;
    251: T0 = 32'hcc57b563;
    252: T0 = 32'hcdcf097d;
    253: T0 = 32'ha0f782ac;
    254: T0 = 32'h229168b7;
    255: T0 = 32'h689f7cde;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[7:0];
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T6 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_32(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[7:0] T5;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T6;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (T5)
    0: T0 = 32'hdca1ecb1;
    1: T0 = 32'h61b28272;
    2: T0 = 32'hb6a1a44a;
    3: T0 = 32'h92bb4688;
    4: T0 = 32'h36b8daf1;
    5: T0 = 32'hface272c;
    6: T0 = 32'h51ddfe4d;
    7: T0 = 32'h436c0f5;
    8: T0 = 32'h39a73450;
    9: T0 = 32'h4644d473;
    10: T0 = 32'h540c3900;
    11: T0 = 32'he06b0e2e;
    12: T0 = 32'hb464fb89;
    13: T0 = 32'hd3615f7;
    14: T0 = 32'hd25fd3d8;
    15: T0 = 32'h75e121a2;
    16: T0 = 32'h375e61bb;
    17: T0 = 32'h619b13aa;
    18: T0 = 32'ha782b6f0;
    19: T0 = 32'h82c20a6c;
    20: T0 = 32'hb7fc8ae1;
    21: T0 = 32'hd2c57dee;
    22: T0 = 32'h19e4e666;
    23: T0 = 32'he56eb9ac;
    24: T0 = 32'hb1f093d0;
    25: T0 = 32'hbe40f30b;
    26: T0 = 32'h23cee2f3;
    27: T0 = 32'ha26b3026;
    28: T0 = 32'ha2669188;
    29: T0 = 32'h2aa9d75f;
    30: T0 = 32'he64f2561;
    31: T0 = 32'hc1d56d66;
    32: T0 = 32'hc56f8e40;
    33: T0 = 32'h7be89343;
    34: T0 = 32'h7d75cc3d;
    35: T0 = 32'h1aaba413;
    36: T0 = 32'h9cf3b251;
    37: T0 = 32'h2b1a3544;
    38: T0 = 32'h5fdad955;
    39: T0 = 32'h30760a83;
    40: T0 = 32'h6e8756d6;
    41: T0 = 32'hc60684a2;
    42: T0 = 32'h151f7d64;
    43: T0 = 32'hc47d8649;
    44: T0 = 32'h3c60bf98;
    45: T0 = 32'h597509b4;
    46: T0 = 32'hd2aedb28;
    47: T0 = 32'h7121f627;
    48: T0 = 32'hface11af;
    49: T0 = 32'h5ec26edc;
    50: T0 = 32'hda796545;
    51: T0 = 32'h9aba912f;
    52: T0 = 32'hecd30dee;
    53: T0 = 32'h7ab1c30b;
    54: T0 = 32'h1ffc2fc9;
    55: T0 = 32'h9276e97c;
    56: T0 = 32'h3e8b89a1;
    57: T0 = 32'h56563e79;
    58: T0 = 32'hc2174392;
    59: T0 = 32'hfc2d61bc;
    60: T0 = 32'hbb3100e7;
    61: T0 = 32'h5feedd89;
    62: T0 = 32'hd7fbb25e;
    63: T0 = 32'h35a10931;
    64: T0 = 32'hbfdefeb0;
    65: T0 = 32'h5c3bc47;
    66: T0 = 32'he2f91ab1;
    67: T0 = 32'he03eb516;
    68: T0 = 32'h42b8b15a;
    69: T0 = 32'hbef59c7a;
    70: T0 = 32'h5f2dd900;
    71: T0 = 32'h80bf1d9e;
    72: T0 = 32'h7203cf9f;
    73: T0 = 32'h54f67caa;
    74: T0 = 32'hc20ccd56;
    75: T0 = 32'h39a99265;
    76: T0 = 32'h1db1e510;
    77: T0 = 32'h1daeb8d3;
    78: T0 = 32'hcfff49ad;
    79: T0 = 32'hbdc94625;
    80: T0 = 32'h239a68f3;
    81: T0 = 32'h2c4992a2;
    82: T0 = 32'h94308f42;
    83: T0 = 32'ha94766f0;
    84: T0 = 32'h6e1152c5;
    85: T0 = 32'h586fade4;
    86: T0 = 32'h27a5c76e;
    87: T0 = 32'hb55c72f9;
    88: T0 = 32'h63411cf8;
    89: T0 = 32'h34f7c1d4;
    90: T0 = 32'hb1cea20d;
    91: T0 = 32'h212e5a64;
    92: T0 = 32'h8dc13f88;
    93: T0 = 32'h4f3fae7c;
    94: T0 = 32'h4e3cc8d1;
    95: T0 = 32'hfa1a8582;
    96: T0 = 32'hb19a7bd0;
    97: T0 = 32'heae33404;
    98: T0 = 32'h26f822a3;
    99: T0 = 32'h87cbb73c;
    100: T0 = 32'h5e8c814a;
    101: T0 = 32'hcc3fd8fb;
    102: T0 = 32'h26131509;
    103: T0 = 32'haad8afd2;
    104: T0 = 32'hd7748a2d;
    105: T0 = 32'hf0723dca;
    106: T0 = 32'hdb318956;
    107: T0 = 32'h1f988ce7;
    108: T0 = 32'h4db24c17;
    109: T0 = 32'h49471299;
    110: T0 = 32'h546a489e;
    111: T0 = 32'hf6d8425c;
    112: T0 = 32'h29d8f9a8;
    113: T0 = 32'h17441f46;
    114: T0 = 32'h64f53ac1;
    115: T0 = 32'h493f9f27;
    116: T0 = 32'h69638300;
    117: T0 = 32'h65bfadc2;
    118: T0 = 32'hd203777b;
    119: T0 = 32'h18b38acc;
    120: T0 = 32'h6e1bcb8f;
    121: T0 = 32'h402fe5b6;
    122: T0 = 32'hbdd0055;
    123: T0 = 32'h5fae2262;
    124: T0 = 32'hfd993250;
    125: T0 = 32'h7c77b38c;
    126: T0 = 32'h88b14b55;
    127: T0 = 32'h1ebed465;
    128: T0 = 32'h7b98eef1;
    129: T0 = 32'hecc85652;
    130: T0 = 32'ha13e8840;
    131: T0 = 32'h3f431e03;
    132: T0 = 32'h9710c801;
    133: T0 = 32'hb1483d40;
    134: T0 = 32'hefa49a77;
    135: T0 = 32'hf748049d;
    136: T0 = 32'hd9e05f5e;
    137: T0 = 32'hb8814476;
    138: T0 = 32'hb48a684d;
    139: T0 = 32'h51002265;
    140: T0 = 32'h8c427788;
    141: T0 = 32'h8131b9a4;
    142: T0 = 32'h66c651e9;
    143: T0 = 32'hfb4ef424;
    144: T0 = 32'he0e3de11;
    145: T0 = 32'heef3186d;
    146: T0 = 32'h9e524c38;
    147: T0 = 32'h8c88bd53;
    148: T0 = 32'hbe134150;
    149: T0 = 32'hc8059c7c;
    150: T0 = 32'h25c2d017;
    151: T0 = 32'hde758d9f;
    152: T0 = 32'h6ddcf1f;
    153: T0 = 32'h5fdec8e2;
    154: T0 = 32'h44729d5c;
    155: T0 = 32'he84c9a65;
    156: T0 = 32'h267e788;
    157: T0 = 32'h77892811;
    158: T0 = 32'hb9bc48af;
    159: T0 = 32'h52a1d6a4;
    160: T0 = 32'hf50668e8;
    161: T0 = 32'h33be1972;
    162: T0 = 32'h6ec41bc1;
    163: T0 = 32'h23e0df76;
    164: T0 = 32'h90ee0101;
    165: T0 = 32'h8d8eade2;
    166: T0 = 32'hc01bf76e;
    167: T0 = 32'h26abbae4;
    168: T0 = 32'hac7cab15;
    169: T0 = 32'h8b297137;
    170: T0 = 32'h7b59a045;
    171: T0 = 32'hc7d22242;
    172: T0 = 32'h41bc9271;
    173: T0 = 32'h64c7a2ac;
    174: T0 = 32'hb7c96111;
    175: T0 = 32'h2dcdce4;
    176: T0 = 32'he585ff1;
    177: T0 = 32'h11b79ce6;
    178: T0 = 32'h6e884ae2;
    179: T0 = 32'h7709733;
    180: T0 = 32'ha3ee904e;
    181: T0 = 32'h8ece00fc;
    182: T0 = 32'h505a1714;
    183: T0 = 32'h22a32791;
    184: T0 = 32'hb13e668f;
    185: T0 = 32'h8f893cca;
    186: T0 = 32'h474ce146;
    187: T0 = 32'hc3f22f66;
    188: T0 = 32'h51346d4f;
    189: T0 = 32'h24c612a9;
    190: T0 = 32'hb35b78f6;
    191: T0 = 32'h4ccf45e;
    192: T0 = 32'hf55934e;
    193: T0 = 32'h926f5d4f;
    194: T0 = 32'h4fd97db5;
    195: T0 = 32'h4d1e9127;
    196: T0 = 32'h418fa70a;
    197: T0 = 32'hce3cf22b;
    198: T0 = 32'h35137191;
    199: T0 = 32'haad9492a;
    200: T0 = 32'h65d89af;
    201: T0 = 32'h7d3e7eb8;
    202: T0 = 32'h46315f96;
    203: T0 = 32'h77a8c8ca;
    204: T0 = 32'h5b1a8070;
    205: T0 = 32'h7247ef81;
    206: T0 = 32'h1d84262e;
    207: T0 = 32'h16bac6a1;
    208: T0 = 32'hbb9885bd;
    209: T0 = 32'h9607aa82;
    210: T0 = 32'h7e59e544;
    211: T0 = 32'h4c3db328;
    212: T0 = 32'h601b9ce4;
    213: T0 = 32'hefb12164;
    214: T0 = 32'hde1d47cd;
    215: T0 = 32'hd89581f9;
    216: T0 = 32'h4d1f3fc9;
    217: T0 = 32'h465f2648;
    218: T0 = 32'hce2263e0;
    219: T0 = 32'h5fbe422e;
    220: T0 = 32'h9b99b3a9;
    221: T0 = 32'hf58eef9e;
    222: T0 = 32'ha973b7c4;
    223: T0 = 32'h178a0427;
    224: T0 = 32'h3ba1eac3;
    225: T0 = 32'h7fe8c4b0;
    226: T0 = 32'hcc2583c2;
    227: T0 = 32'h1ac35ddc;
    228: T0 = 32'hbdf348ef;
    229: T0 = 32'h71480e93;
    230: T0 = 32'h89e4ae6a;
    231: T0 = 32'h153ed7d0;
    232: T0 = 32'h2fc1703b;
    233: T0 = 32'h6a874947;
    234: T0 = 32'ha18ea40d;
    235: T0 = 32'h846f7f93;
    236: T0 = 32'ha7626cc7;
    237: T0 = 32'h1d7b1478;
    238: T0 = 32'h42a8c8b7;
    239: T0 = 32'h681729d8;
    240: T0 = 32'hfcdecce9;
    241: T0 = 32'hda480376;
    242: T0 = 32'h1cb68cc7;
    243: T0 = 32'h4d445c01;
    244: T0 = 32'hfd476805;
    245: T0 = 32'h4520a700;
    246: T0 = 32'hac73fa5c;
    247: T0 = 32'hdf4ac2c1;
    248: T0 = 32'h865c7876;
    249: T0 = 32'hd93d4433;
    250: T0 = 32'h6bf1a60d;
    251: T0 = 32'he542f12;
    252: T0 = 32'h9b4b7b79;
    253: T0 = 32'he2c1192c;
    254: T0 = 32'hbc00f410;
    255: T0 = 32'hcabfb8a2;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[7:0];
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T6 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_33(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[7:0] T5;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T6;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (T5)
    0: T0 = 32'h239a86cf;
    1: T0 = 32'h170643fb;
    2: T0 = 32'h78cdbc0e;
    3: T0 = 32'h643c40c3;
    4: T0 = 32'h61e22eb5;
    5: T0 = 32'h27b12d24;
    6: T0 = 32'hd80deaf7;
    7: T0 = 32'h49b7c2a9;
    8: T0 = 32'h4a2b5550;
    9: T0 = 32'h11e95335;
    10: T0 = 32'hcbdc3aa9;
    11: T0 = 32'h7faa521a;
    12: T0 = 32'hd1999b98;
    13: T0 = 32'hb4be8d66;
    14: T0 = 32'hadb2a761;
    15: T0 = 32'h60ea9a2;
    16: T0 = 32'hf83f1b7;
    17: T0 = 32'h7fea6c85;
    18: T0 = 32'hfd4022b0;
    19: T0 = 32'h3ae136ae;
    20: T0 = 32'h36b288de;
    21: T0 = 32'hb10a515a;
    22: T0 = 32'h59cc2ea2;
    23: T0 = 32'h153e15be;
    24: T0 = 32'hfbc7868c;
    25: T0 = 32'h4ec74769;
    26: T0 = 32'h948fc3fb;
    27: T0 = 32'hc4656124;
    28: T0 = 32'ha4606cc6;
    29: T0 = 32'h1836915b;
    30: T0 = 32'h42ce11fe;
    31: T0 = 32'h79452f5c;
    32: T0 = 32'hd6ccb0af;
    33: T0 = 32'h61bfabbb;
    34: T0 = 32'h6cb8270f;
    35: T0 = 32'h13e28a4e;
    36: T0 = 32'h19fead2e;
    37: T0 = 32'h45aeee23;
    38: T0 = 32'hca8b6eeb;
    39: T0 = 32'h26aad560;
    40: T0 = 32'hf77cb9b1;
    41: T0 = 32'ha9217f29;
    42: T0 = 32'h5b4dd392;
    43: T0 = 32'h82db4d9a;
    44: T0 = 32'h6992c151;
    45: T0 = 32'h44f3754a;
    46: T0 = 32'hd74ab458;
    47: T0 = 32'ha45708f0;
    48: T0 = 32'h8850ee68;
    49: T0 = 32'h722e5e52;
    50: T0 = 32'h4dbf3844;
    51: T0 = 32'h13893c17;
    52: T0 = 32'h89cec804;
    53: T0 = 32'h678e25d2;
    54: T0 = 32'head3be74;
    55: T0 = 32'h667a0ad5;
    56: T0 = 32'hbf4cefde;
    57: T0 = 32'h892f24f3;
    58: T0 = 32'h7b112c55;
    59: T0 = 32'h9e9b0362;
    60: T0 = 32'h79927ac9;
    61: T0 = 32'hd05119a4;
    62: T0 = 32'hf74adab1;
    63: T0 = 32'h2431f50c;
    64: T0 = 32'hc8e0fcc8;
    65: T0 = 32'hfac1b13f;
    66: T0 = 32'h203d3abf;
    67: T0 = 32'h8fab9e11;
    68: T0 = 32'h4c0cb350;
    69: T0 = 32'hb8f37f2c;
    70: T0 = 32'hdebdd915;
    71: T0 = 32'hba91cb83;
    72: T0 = 32'hc72756d3;
    73: T0 = 32'h7433f4aa;
    74: T0 = 32'hdda3e925;
    75: T0 = 32'hde039063;
    76: T0 = 32'h5d928b38;
    77: T0 = 32'hcd4763e6;
    78: T0 = 32'h54737968;
    79: T0 = 32'hfc9a62e7;
    80: T0 = 32'h39d2c8ba;
    81: T0 = 32'h1f461f42;
    82: T0 = 32'h7cc5f8d0;
    83: T0 = 32'h4838b757;
    84: T0 = 32'h6cf39a40;
    85: T0 = 32'h579f39e0;
    86: T0 = 32'h505fd7ee;
    87: T0 = 32'h10b798bd;
    88: T0 = 32'hf1b8bcc;
    89: T0 = 32'h47ef647a;
    90: T0 = 32'h4a0ce275;
    91: T0 = 32'h5decb266;
    92: T0 = 32'hf3b5b218;
    93: T0 = 32'hbcaea3ce;
    94: T0 = 32'h89314561;
    95: T0 = 32'h1ca7d627;
    96: T0 = 32'h179fd891;
    97: T0 = 32'h31eef405;
    98: T0 = 32'hbfacc6c;
    99: T0 = 32'h1bc17754;
    100: T0 = 32'h9976d0da;
    101: T0 = 32'h2f859af9;
    102: T0 = 32'h2d821101;
    103: T0 = 32'hf67a151a;
    104: T0 = 32'h7acc070d;
    105: T0 = 32'h6916a8e2;
    106: T0 = 32'h531da94e;
    107: T0 = 32'h82b9cded;
    108: T0 = 32'h7272e58e;
    109: T0 = 32'h1070aa31;
    110: T0 = 32'hd53ec8be;
    111: T0 = 32'h2551071e;
    112: T0 = 32'hfce013e6;
    113: T0 = 32'h61b06cc5;
    114: T0 = 32'h96825bb3;
    115: T0 = 32'ha040b9b7;
    116: T0 = 32'hb72a258a;
    117: T0 = 32'h8ac6d15b;
    118: T0 = 32'h39e21493;
    119: T0 = 32'h47882f06;
    120: T0 = 32'h39f8ca2f;
    121: T0 = 32'h8788438e;
    122: T0 = 32'h26c8cf7e;
    123: T0 = 32'he271e5d1;
    124: T0 = 32'h62642476;
    125: T0 = 32'h2689928f;
    126: T0 = 32'hbbce283f;
    127: T0 = 32'hc3c45e1c;
    128: T0 = 32'h4645feb0;
    129: T0 = 32'h7ee9d47;
    130: T0 = 32'he5d518b9;
    131: T0 = 32'hb3afb516;
    132: T0 = 32'h12b9a15a;
    133: T0 = 32'hbe5f9c78;
    134: T0 = 32'h538dd800;
    135: T0 = 32'h3ebc9d9f;
    136: T0 = 32'hfb43cf9d;
    137: T0 = 32'h64a22ca2;
    138: T0 = 32'h948fcc66;
    139: T0 = 32'he62e8241;
    140: T0 = 32'h2da0e5c0;
    141: T0 = 32'hd7f31db;
    142: T0 = 32'h42cf49a4;
    143: T0 = 32'h795e4665;
    144: T0 = 32'h3b5a3322;
    145: T0 = 32'h3f46adad;
    146: T0 = 32'h65f113b1;
    147: T0 = 32'h1bb389fe;
    148: T0 = 32'h78f1e5ee;
    149: T0 = 32'h7795dabb;
    150: T0 = 32'h5e890522;
    151: T0 = 32'h95767f2a;
    152: T0 = 32'h6e03a0a3;
    153: T0 = 32'h646ebbcc;
    154: T0 = 32'h819d8ebb;
    155: T0 = 32'ha42dddf0;
    156: T0 = 32'hbdf10cf6;
    157: T0 = 32'h5e3fe65b;
    158: T0 = 32'h822c283f;
    159: T0 = 32'hd9030ad8;
    160: T0 = 32'hfbda9c15;
    161: T0 = 32'hb1b6f00d;
    162: T0 = 32'h7a8bec2c;
    163: T0 = 32'h21707608;
    164: T0 = 32'h13eed07b;
    165: T0 = 32'h8cfe9259;
    166: T0 = 32'h51da0981;
    167: T0 = 32'h66a20533;
    168: T0 = 32'h3d3e96e9;
    169: T0 = 32'h87a9ace0;
    170: T0 = 32'h424c7946;
    171: T0 = 32'hcbda8dcd;
    172: T0 = 32'h71bced8f;
    173: T0 = 32'h24c20cb1;
    174: T0 = 32'hb5dfdabe;
    175: T0 = 32'h6e5231b;
    176: T0 = 32'h75d1c6c;
    177: T0 = 32'h154e55d4;
    178: T0 = 32'hf389e847;
    179: T0 = 32'hd93f6481;
    180: T0 = 32'h60f11505;
    181: T0 = 32'h76b5a105;
    182: T0 = 32'he92d1bdd;
    183: T0 = 32'h91ff4a41;
    184: T0 = 32'h6a236c6e;
    185: T0 = 32'h14ea04bf;
    186: T0 = 32'hc39c6504;
    187: T0 = 32'h36a96799;
    188: T0 = 32'hd0d93abf;
    189: T0 = 32'hbbbe08a4;
    190: T0 = 32'hcf769a1e;
    191: T0 = 32'h8741f49f;
    192: T0 = 32'h298bd606;
    193: T0 = 32'hec997859;
    194: T0 = 32'hb1274c3d;
    195: T0 = 32'haead200b;
    196: T0 = 32'h9610b7b1;
    197: T0 = 32'hba5ade5d;
    198: T0 = 32'h13bcd895;
    199: T0 = 32'hfc04061e;
    200: T0 = 32'hd1a6477e;
    201: T0 = 32'h3491cc27;
    202: T0 = 32'hb4a25ff8;
    203: T0 = 32'h7924d399;
    204: T0 = 32'h806ef51e;
    205: T0 = 32'hcd185db1;
    206: T0 = 32'h56f717ea;
    207: T0 = 32'hfb6813b1;
    208: T0 = 32'h2363de49;
    209: T0 = 32'hf8b3f955;
    210: T0 = 32'h180e6c0f;
    211: T0 = 32'h2740ed01;
    212: T0 = 32'h9f0e0138;
    213: T0 = 32'h80eaa615;
    214: T0 = 32'h9472d951;
    215: T0 = 32'h6f02ce05;
    216: T0 = 32'h95bc49bf;
    217: T0 = 32'h9b998ce3;
    218: T0 = 32'hf4685d14;
    219: T0 = 32'hcb538fdb;
    220: T0 = 32'h266e911;
    221: T0 = 32'he6c03890;
    222: T0 = 32'hf7d3dabe;
    223: T0 = 32'h64fcf8b0;
    224: T0 = 32'hc465de51;
    225: T0 = 32'h6fb2dc07;
    226: T0 = 32'h9f434820;
    227: T0 = 32'h1ab97d73;
    228: T0 = 32'h1ed351db;
    229: T0 = 32'hfb5a985a;
    230: T0 = 32'h5dfc9135;
    231: T0 = 32'h9032071f;
    232: T0 = 32'h3f8f47ef;
    233: T0 = 32'h464689e4;
    234: T0 = 32'h702f8d5d;
    235: T0 = 32'hcc6fbbf9;
    236: T0 = 32'hb060a68e;
    237: T0 = 32'h155eaab1;
    238: T0 = 32'hd1e748ae;
    239: T0 = 32'h6561569f;
    240: T0 = 32'h774e0dce;
    241: T0 = 32'h64767e5;
    242: T0 = 32'he0b9bbaf;
    243: T0 = 32'hc53a16b8;
    244: T0 = 32'h6ad8be5e;
    245: T0 = 32'h7eff539d;
    246: T0 = 32'h523d24d8;
    247: T0 = 32'h20c5efc3;
    248: T0 = 32'h553364a6;
    249: T0 = 32'h1430940f;
    250: T0 = 32'hdb05e12e;
    251: T0 = 32'h37aa65f0;
    252: T0 = 32'hdd990936;
    253: T0 = 32'hcfee50cf;
    254: T0 = 32'h4c73b95e;
    255: T0 = 32'h95aa23da;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[7:0];
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T6 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_34(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[7:0] io_weights
);

  reg [7:0] weightsReg;
  wire[7:0] T4;
  reg [7:0] T0;
  wire[7:0] T5;
  wire[8:0] addr;
  reg [8:0] counter;
  wire[8:0] T6;
  wire[8:0] T2;
  wire[8:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 8'h0 : T0;
  always @(*) case (T5)
    0: T0 = 8'hb;
    1: T0 = 8'hf4;
    2: T0 = 8'hf5;
    3: T0 = 8'h7;
    4: T0 = 8'hfa;
    5: T0 = 8'ha;
    6: T0 = 8'hff;
    7: T0 = 8'hfc;
    8: T0 = 8'h1;
    9: T0 = 8'h2;
    10: T0 = 8'hfb;
    11: T0 = 8'h0;
    12: T0 = 8'h3;
    13: T0 = 8'h2;
    14: T0 = 8'hc;
    15: T0 = 8'h2;
    16: T0 = 8'h1;
    17: T0 = 8'h4;
    18: T0 = 8'h0;
    19: T0 = 8'h3;
    20: T0 = 8'hfb;
    21: T0 = 8'hf8;
    22: T0 = 8'hfe;
    23: T0 = 8'hf0;
    24: T0 = 8'hc;
    25: T0 = 8'hf9;
    26: T0 = 8'hfa;
    27: T0 = 8'hfe;
    28: T0 = 8'h10;
    29: T0 = 8'h8;
    30: T0 = 8'hfd;
    31: T0 = 8'hff;
    32: T0 = 8'h7;
    33: T0 = 8'hfc;
    34: T0 = 8'h3;
    35: T0 = 8'h5;
    36: T0 = 8'h9;
    37: T0 = 8'h2;
    38: T0 = 8'h0;
    39: T0 = 8'hf4;
    40: T0 = 8'hfa;
    41: T0 = 8'hf7;
    42: T0 = 8'h4;
    43: T0 = 8'h6;
    44: T0 = 8'h3;
    45: T0 = 8'hf9;
    46: T0 = 8'hfb;
    47: T0 = 8'hfc;
    48: T0 = 8'hfe;
    49: T0 = 8'hf6;
    50: T0 = 8'h1;
    51: T0 = 8'hfe;
    52: T0 = 8'h3f;
    53: T0 = 8'h6;
    54: T0 = 8'h1;
    55: T0 = 8'hf7;
    56: T0 = 8'h3;
    57: T0 = 8'h1;
    58: T0 = 8'hf4;
    59: T0 = 8'h3;
    60: T0 = 8'hf8;
    61: T0 = 8'h6;
    62: T0 = 8'h1;
    63: T0 = 8'hf8;
    64: T0 = 8'hfd;
    65: T0 = 8'hf9;
    66: T0 = 8'h6;
    67: T0 = 8'hf8;
    68: T0 = 8'h1;
    69: T0 = 8'hf6;
    70: T0 = 8'ha;
    71: T0 = 8'hf8;
    72: T0 = 8'hff;
    73: T0 = 8'hd;
    74: T0 = 8'hfa;
    75: T0 = 8'hfc;
    76: T0 = 8'hf6;
    77: T0 = 8'h8;
    78: T0 = 8'hf3;
    79: T0 = 8'h5;
    80: T0 = 8'hff;
    81: T0 = 8'hff;
    82: T0 = 8'hfe;
    83: T0 = 8'hf3;
    84: T0 = 8'h2;
    85: T0 = 8'h3;
    86: T0 = 8'hff;
    87: T0 = 8'hf9;
    88: T0 = 8'h4;
    89: T0 = 8'h7;
    90: T0 = 8'hf9;
    91: T0 = 8'hff;
    92: T0 = 8'h6;
    93: T0 = 8'hfd;
    94: T0 = 8'h2;
    95: T0 = 8'h4;
    96: T0 = 8'h12;
    97: T0 = 8'hff;
    98: T0 = 8'h2;
    99: T0 = 8'hff;
    100: T0 = 8'hfc;
    101: T0 = 8'h0;
    102: T0 = 8'h1;
    103: T0 = 8'hf9;
    104: T0 = 8'hd;
    105: T0 = 8'hd;
    106: T0 = 8'hfb;
    107: T0 = 8'h11;
    108: T0 = 8'hf6;
    109: T0 = 8'hfc;
    110: T0 = 8'h2;
    111: T0 = 8'h0;
    112: T0 = 8'hff;
    113: T0 = 8'h2;
    114: T0 = 8'h0;
    115: T0 = 8'hfc;
    116: T0 = 8'hff;
    117: T0 = 8'hfd;
    118: T0 = 8'h3;
    119: T0 = 8'hf8;
    120: T0 = 8'hfc;
    121: T0 = 8'hf3;
    122: T0 = 8'hfc;
    123: T0 = 8'hfd;
    124: T0 = 8'hf9;
    125: T0 = 8'hfa;
    126: T0 = 8'hf8;
    127: T0 = 8'hfe;
    128: T0 = 8'h4;
    129: T0 = 8'hff;
    130: T0 = 8'h8;
    131: T0 = 8'h2;
    132: T0 = 8'h9;
    133: T0 = 8'h4;
    134: T0 = 8'h0;
    135: T0 = 8'hf9;
    136: T0 = 8'hf8;
    137: T0 = 8'h1;
    138: T0 = 8'h2;
    139: T0 = 8'hfb;
    140: T0 = 8'h4;
    141: T0 = 8'hfe;
    142: T0 = 8'hf9;
    143: T0 = 8'hfd;
    144: T0 = 8'hfb;
    145: T0 = 8'hc;
    146: T0 = 8'h4;
    147: T0 = 8'hf9;
    148: T0 = 8'h7;
    149: T0 = 8'hfb;
    150: T0 = 8'hfb;
    151: T0 = 8'h3;
    152: T0 = 8'hfc;
    153: T0 = 8'h1;
    154: T0 = 8'h2;
    155: T0 = 8'hfd;
    156: T0 = 8'h2;
    157: T0 = 8'h6;
    158: T0 = 8'hfb;
    159: T0 = 8'hff;
    160: T0 = 8'hfc;
    161: T0 = 8'h3;
    162: T0 = 8'hfd;
    163: T0 = 8'hf8;
    164: T0 = 8'ha;
    165: T0 = 8'hfc;
    166: T0 = 8'hfd;
    167: T0 = 8'h2;
    168: T0 = 8'h8;
    169: T0 = 8'h5;
    170: T0 = 8'hfa;
    171: T0 = 8'h6;
    172: T0 = 8'h0;
    173: T0 = 8'hfb;
    174: T0 = 8'hfe;
    175: T0 = 8'h0;
    176: T0 = 8'h5;
    177: T0 = 8'hee;
    178: T0 = 8'hfa;
    179: T0 = 8'hff;
    180: T0 = 8'h4;
    181: T0 = 8'hfb;
    182: T0 = 8'h8;
    183: T0 = 8'hf5;
    184: T0 = 8'ha;
    185: T0 = 8'h7;
    186: T0 = 8'h6;
    187: T0 = 8'h4;
    188: T0 = 8'hfe;
    189: T0 = 8'h2;
    190: T0 = 8'hf4;
    191: T0 = 8'h7;
    192: T0 = 8'h5;
    193: T0 = 8'h9;
    194: T0 = 8'h0;
    195: T0 = 8'h1;
    196: T0 = 8'hfe;
    197: T0 = 8'hf9;
    198: T0 = 8'hfd;
    199: T0 = 8'hfc;
    200: T0 = 8'hff;
    201: T0 = 8'h4;
    202: T0 = 8'h9;
    203: T0 = 8'hf7;
    204: T0 = 8'hf7;
    205: T0 = 8'hfc;
    206: T0 = 8'h1;
    207: T0 = 8'hfa;
    208: T0 = 8'hfe;
    209: T0 = 8'hfc;
    210: T0 = 8'hfb;
    211: T0 = 8'h4;
    212: T0 = 8'h1;
    213: T0 = 8'hff;
    214: T0 = 8'h1;
    215: T0 = 8'hc;
    216: T0 = 8'h3;
    217: T0 = 8'hff;
    218: T0 = 8'hf4;
    219: T0 = 8'h8;
    220: T0 = 8'h3;
    221: T0 = 8'h3;
    222: T0 = 8'hf6;
    223: T0 = 8'hff;
    224: T0 = 8'h8;
    225: T0 = 8'h6;
    226: T0 = 8'h1;
    227: T0 = 8'h6;
    228: T0 = 8'h1;
    229: T0 = 8'h7;
    230: T0 = 8'hfc;
    231: T0 = 8'ha;
    232: T0 = 8'h5;
    233: T0 = 8'h6;
    234: T0 = 8'h3;
    235: T0 = 8'hf4;
    236: T0 = 8'hfd;
    237: T0 = 8'hf2;
    238: T0 = 8'hfe;
    239: T0 = 8'hff;
    240: T0 = 8'hf8;
    241: T0 = 8'hfc;
    242: T0 = 8'h4;
    243: T0 = 8'hfc;
    244: T0 = 8'hf7;
    245: T0 = 8'hfe;
    246: T0 = 8'hfd;
    247: T0 = 8'hf8;
    248: T0 = 8'hf9;
    249: T0 = 8'hfc;
    250: T0 = 8'hf1;
    251: T0 = 8'hfc;
    252: T0 = 8'hfc;
    253: T0 = 8'hff;
    254: T0 = 8'hf8;
    255: T0 = 8'h5;
    default: begin
      T0 = 8'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[7:0];
  assign addr = io_restartIn ? 9'h0 : counter;
  assign T6 = reset ? 9'h0 : T2;
  assign T2 = io_restartIn ? 9'h1 : T3;
  assign T3 = counter + 9'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 8'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 9'h0;
    end else if(io_restartIn) begin
      counter <= 9'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryStreamer_2(input clk, input reset,
    input  io_restart,
    output[15:0] io_weights_15,
    output[15:0] io_weights_14,
    output[15:0] io_weights_13,
    output[15:0] io_weights_12,
    output[15:0] io_weights_11,
    output[15:0] io_weights_10,
    output[15:0] io_weights_9,
    output[15:0] io_weights_8,
    output[15:0] io_weights_7,
    output[15:0] io_weights_6,
    output[15:0] io_weights_5,
    output[15:0] io_weights_4,
    output[15:0] io_weights_3,
    output[15:0] io_weights_2,
    output[15:0] io_weights_1,
    output[15:0] io_weights_0,
    output[7:0] io_bias
);

  wire[7:0] T18;
  wire[8:0] T0;
  wire[8:0] T1;
  wire[15:0] T2;
  wire[15:0] T3;
  wire[15:0] T4;
  wire[15:0] T5;
  wire[15:0] T6;
  wire[15:0] T7;
  wire[15:0] T8;
  wire[15:0] T9;
  wire[15:0] T10;
  wire[15:0] T11;
  wire[15:0] T12;
  wire[15:0] T13;
  wire[15:0] T14;
  wire[15:0] T15;
  wire[15:0] T16;
  wire[15:0] T17;
  wire MemoryUnit_io_restartOut;
  wire[31:0] MemoryUnit_io_weights;
  wire MemoryUnit_1_io_restartOut;
  wire[31:0] MemoryUnit_1_io_weights;
  wire MemoryUnit_2_io_restartOut;
  wire[31:0] MemoryUnit_2_io_weights;
  wire MemoryUnit_3_io_restartOut;
  wire[31:0] MemoryUnit_3_io_weights;
  wire MemoryUnit_4_io_restartOut;
  wire[31:0] MemoryUnit_4_io_weights;
  wire MemoryUnit_5_io_restartOut;
  wire[31:0] MemoryUnit_5_io_weights;
  wire MemoryUnit_6_io_restartOut;
  wire[31:0] MemoryUnit_6_io_weights;
  wire[31:0] MemoryUnit_7_io_weights;
  wire[7:0] biasMemoryUnit_io_weights;


  assign io_bias = T18;
  assign T18 = T0[7:0];
  assign T0 = T1;
  assign T1 = {1'h0, biasMemoryUnit_io_weights};
  assign io_weights_0 = T2;
  assign T2 = MemoryUnit_io_weights[15:0];
  assign io_weights_1 = T3;
  assign T3 = MemoryUnit_io_weights[31:16];
  assign io_weights_2 = T4;
  assign T4 = MemoryUnit_1_io_weights[15:0];
  assign io_weights_3 = T5;
  assign T5 = MemoryUnit_1_io_weights[31:16];
  assign io_weights_4 = T6;
  assign T6 = MemoryUnit_2_io_weights[15:0];
  assign io_weights_5 = T7;
  assign T7 = MemoryUnit_2_io_weights[31:16];
  assign io_weights_6 = T8;
  assign T8 = MemoryUnit_3_io_weights[15:0];
  assign io_weights_7 = T9;
  assign T9 = MemoryUnit_3_io_weights[31:16];
  assign io_weights_8 = T10;
  assign T10 = MemoryUnit_4_io_weights[15:0];
  assign io_weights_9 = T11;
  assign T11 = MemoryUnit_4_io_weights[31:16];
  assign io_weights_10 = T12;
  assign T12 = MemoryUnit_5_io_weights[15:0];
  assign io_weights_11 = T13;
  assign T13 = MemoryUnit_5_io_weights[31:16];
  assign io_weights_12 = T14;
  assign T14 = MemoryUnit_6_io_weights[15:0];
  assign io_weights_13 = T15;
  assign T15 = MemoryUnit_6_io_weights[31:16];
  assign io_weights_14 = T16;
  assign T16 = MemoryUnit_7_io_weights[15:0];
  assign io_weights_15 = T17;
  assign T17 = MemoryUnit_7_io_weights[31:16];
  MemoryUnit_26 MemoryUnit(.clk(clk), .reset(reset),
       .io_restartIn( io_restart ),
       .io_restartOut( MemoryUnit_io_restartOut ),
       .io_weights( MemoryUnit_io_weights )
  );
  MemoryUnit_27 MemoryUnit_1(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_io_restartOut ),
       .io_restartOut( MemoryUnit_1_io_restartOut ),
       .io_weights( MemoryUnit_1_io_weights )
  );
  MemoryUnit_28 MemoryUnit_2(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_1_io_restartOut ),
       .io_restartOut( MemoryUnit_2_io_restartOut ),
       .io_weights( MemoryUnit_2_io_weights )
  );
  MemoryUnit_29 MemoryUnit_3(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_2_io_restartOut ),
       .io_restartOut( MemoryUnit_3_io_restartOut ),
       .io_weights( MemoryUnit_3_io_weights )
  );
  MemoryUnit_30 MemoryUnit_4(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_3_io_restartOut ),
       .io_restartOut( MemoryUnit_4_io_restartOut ),
       .io_weights( MemoryUnit_4_io_weights )
  );
  MemoryUnit_31 MemoryUnit_5(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_4_io_restartOut ),
       .io_restartOut( MemoryUnit_5_io_restartOut ),
       .io_weights( MemoryUnit_5_io_weights )
  );
  MemoryUnit_32 MemoryUnit_6(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_5_io_restartOut ),
       .io_restartOut( MemoryUnit_6_io_restartOut ),
       .io_weights( MemoryUnit_6_io_weights )
  );
  MemoryUnit_33 MemoryUnit_7(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_6_io_restartOut ),
       //.io_restartOut(  )
       .io_weights( MemoryUnit_7_io_weights )
  );
  MemoryUnit_34 biasMemoryUnit(.clk(clk), .reset(reset),
       .io_restartIn( io_restart ),
       //.io_restartOut(  )
       .io_weights( biasMemoryUnit_io_weights )
  );
endmodule

module Warp_2(input clk, input reset,
    input [15:0] io_xIn_2,
    input [15:0] io_xIn_1,
    input [15:0] io_xIn_0,
    input  io_start,
    output io_ready,
    output io_startOut,
    output io_xOut_2,
    output io_xOut_1,
    output io_xOut_0,
    output io_xOutValid,
    input  io_pipeReady,
    output io_done
);

  wire[9:0] T189;
  wire[10:0] T0;
  wire[10:0] T1;
  wire[9:0] T190;
  wire[10:0] T2;
  wire[10:0] T3;
  wire[9:0] T191;
  wire[10:0] T4;
  wire[10:0] T5;
  wire[9:0] T192;
  wire[10:0] T6;
  wire[10:0] T7;
  wire[9:0] T193;
  wire[10:0] T8;
  wire[10:0] T9;
  wire[9:0] T194;
  wire[10:0] T10;
  wire[10:0] T11;
  wire[9:0] T195;
  wire[10:0] T12;
  wire[10:0] T13;
  wire[9:0] T196;
  wire[10:0] T14;
  wire[10:0] T15;
  wire[9:0] T197;
  wire[10:0] T16;
  wire[10:0] T17;
  wire[9:0] T198;
  wire[10:0] T18;
  wire[10:0] T19;
  wire[9:0] T199;
  wire[10:0] T20;
  wire[10:0] T21;
  wire[9:0] T200;
  wire[10:0] T22;
  wire[10:0] T23;
  wire[9:0] T201;
  wire[10:0] T24;
  wire[10:0] T25;
  wire[9:0] T202;
  wire[10:0] T26;
  wire[10:0] T27;
  wire[9:0] T203;
  wire[10:0] T28;
  wire[10:0] T29;
  wire[9:0] T204;
  wire[10:0] T30;
  wire[10:0] T31;
  wire[9:0] T205;
  wire[10:0] T32;
  wire[10:0] T33;
  wire[9:0] T206;
  wire[10:0] T34;
  wire[10:0] T35;
  wire[9:0] T207;
  wire[10:0] T36;
  wire[10:0] T37;
  wire[9:0] T208;
  wire[10:0] T38;
  wire[10:0] T39;
  wire[9:0] T209;
  wire[10:0] T40;
  wire[10:0] T41;
  wire[9:0] T210;
  wire[10:0] T42;
  wire[10:0] T43;
  wire[9:0] T211;
  wire[10:0] T44;
  wire[10:0] T45;
  wire[9:0] T212;
  wire[10:0] T46;
  wire[10:0] T47;
  wire[9:0] T213;
  wire[10:0] T48;
  wire[10:0] T49;
  wire[9:0] T214;
  wire[10:0] T50;
  wire[10:0] T51;
  wire[9:0] T215;
  wire[10:0] T52;
  wire[10:0] T53;
  wire[9:0] T216;
  wire[10:0] T54;
  wire[10:0] T55;
  wire[9:0] T217;
  wire[10:0] T56;
  wire[10:0] T57;
  wire[9:0] T218;
  wire[10:0] T58;
  wire[10:0] T59;
  wire[9:0] T219;
  wire[10:0] T60;
  wire[10:0] T61;
  wire[9:0] T220;
  wire[10:0] T62;
  wire[10:0] T63;
  wire[9:0] T221;
  wire[10:0] T64;
  wire[10:0] T65;
  wire[9:0] T222;
  wire[10:0] T66;
  wire[10:0] T67;
  wire[9:0] T223;
  wire[10:0] T68;
  wire[10:0] T69;
  wire[9:0] T224;
  wire[10:0] T70;
  wire[10:0] T71;
  wire[9:0] T225;
  wire[10:0] T72;
  wire[10:0] T73;
  wire[9:0] T226;
  wire[10:0] T74;
  wire[10:0] T75;
  wire[9:0] T227;
  wire[10:0] T76;
  wire[10:0] T77;
  wire[9:0] T228;
  wire[10:0] T78;
  wire[10:0] T79;
  wire[9:0] T229;
  wire[10:0] T80;
  wire[10:0] T81;
  wire[9:0] T230;
  wire[10:0] T82;
  wire[10:0] T83;
  wire[9:0] T231;
  wire[10:0] T84;
  wire[10:0] T85;
  wire[9:0] T232;
  wire[10:0] T86;
  wire[10:0] T87;
  wire[9:0] T233;
  wire[10:0] T88;
  wire[10:0] T89;
  wire[9:0] T234;
  wire[10:0] T90;
  wire[10:0] T91;
  wire[9:0] T235;
  wire[10:0] T92;
  wire[10:0] T93;
  wire[9:0] T236;
  wire[10:0] T94;
  wire[10:0] T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire[3:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire[3:0] T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire[3:0] T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire Activation_io_out_15;
  wire Activation_io_out_14;
  wire Activation_io_out_13;
  wire Activation_io_out_12;
  wire Activation_io_out_11;
  wire Activation_io_out_10;
  wire Activation_io_out_9;
  wire Activation_io_out_8;
  wire Activation_io_out_7;
  wire Activation_io_out_6;
  wire Activation_io_out_5;
  wire Activation_io_out_4;
  wire Activation_io_out_3;
  wire Activation_io_out_2;
  wire Activation_io_out_1;
  wire Activation_io_out_0;
  wire Activation_1_io_out_15;
  wire Activation_1_io_out_14;
  wire Activation_1_io_out_13;
  wire Activation_1_io_out_12;
  wire Activation_1_io_out_11;
  wire Activation_1_io_out_10;
  wire Activation_1_io_out_9;
  wire Activation_1_io_out_8;
  wire Activation_1_io_out_7;
  wire Activation_1_io_out_6;
  wire Activation_1_io_out_5;
  wire Activation_1_io_out_4;
  wire Activation_1_io_out_3;
  wire Activation_1_io_out_2;
  wire Activation_1_io_out_1;
  wire Activation_1_io_out_0;
  wire Activation_2_io_out_15;
  wire Activation_2_io_out_14;
  wire Activation_2_io_out_13;
  wire Activation_2_io_out_12;
  wire Activation_2_io_out_11;
  wire Activation_2_io_out_10;
  wire Activation_2_io_out_9;
  wire Activation_2_io_out_8;
  wire Activation_2_io_out_7;
  wire Activation_2_io_out_6;
  wire Activation_2_io_out_5;
  wire Activation_2_io_out_4;
  wire Activation_2_io_out_3;
  wire Activation_2_io_out_2;
  wire Activation_2_io_out_1;
  wire Activation_2_io_out_0;
  wire control_io_ready;
  wire control_io_valid;
  wire control_io_done;
  wire[3:0] control_io_selectX;
  wire control_io_memoryRestart;
  wire control_io_chainRestart;
  wire[9:0] Chain_io_ys_15;
  wire[9:0] Chain_io_ys_14;
  wire[9:0] Chain_io_ys_13;
  wire[9:0] Chain_io_ys_12;
  wire[9:0] Chain_io_ys_11;
  wire[9:0] Chain_io_ys_10;
  wire[9:0] Chain_io_ys_9;
  wire[9:0] Chain_io_ys_8;
  wire[9:0] Chain_io_ys_7;
  wire[9:0] Chain_io_ys_6;
  wire[9:0] Chain_io_ys_5;
  wire[9:0] Chain_io_ys_4;
  wire[9:0] Chain_io_ys_3;
  wire[9:0] Chain_io_ys_2;
  wire[9:0] Chain_io_ys_1;
  wire[9:0] Chain_io_ys_0;
  wire[9:0] Chain_1_io_ys_15;
  wire[9:0] Chain_1_io_ys_14;
  wire[9:0] Chain_1_io_ys_13;
  wire[9:0] Chain_1_io_ys_12;
  wire[9:0] Chain_1_io_ys_11;
  wire[9:0] Chain_1_io_ys_10;
  wire[9:0] Chain_1_io_ys_9;
  wire[9:0] Chain_1_io_ys_8;
  wire[9:0] Chain_1_io_ys_7;
  wire[9:0] Chain_1_io_ys_6;
  wire[9:0] Chain_1_io_ys_5;
  wire[9:0] Chain_1_io_ys_4;
  wire[9:0] Chain_1_io_ys_3;
  wire[9:0] Chain_1_io_ys_2;
  wire[9:0] Chain_1_io_ys_1;
  wire[9:0] Chain_1_io_ys_0;
  wire[9:0] Chain_2_io_ys_15;
  wire[9:0] Chain_2_io_ys_14;
  wire[9:0] Chain_2_io_ys_13;
  wire[9:0] Chain_2_io_ys_12;
  wire[9:0] Chain_2_io_ys_11;
  wire[9:0] Chain_2_io_ys_10;
  wire[9:0] Chain_2_io_ys_9;
  wire[9:0] Chain_2_io_ys_8;
  wire[9:0] Chain_2_io_ys_7;
  wire[9:0] Chain_2_io_ys_6;
  wire[9:0] Chain_2_io_ys_5;
  wire[9:0] Chain_2_io_ys_4;
  wire[9:0] Chain_2_io_ys_3;
  wire[9:0] Chain_2_io_ys_2;
  wire[9:0] Chain_2_io_ys_1;
  wire[9:0] Chain_2_io_ys_0;
  wire[15:0] memoryStreamer_io_weights_15;
  wire[15:0] memoryStreamer_io_weights_14;
  wire[15:0] memoryStreamer_io_weights_13;
  wire[15:0] memoryStreamer_io_weights_12;
  wire[15:0] memoryStreamer_io_weights_11;
  wire[15:0] memoryStreamer_io_weights_10;
  wire[15:0] memoryStreamer_io_weights_9;
  wire[15:0] memoryStreamer_io_weights_8;
  wire[15:0] memoryStreamer_io_weights_7;
  wire[15:0] memoryStreamer_io_weights_6;
  wire[15:0] memoryStreamer_io_weights_5;
  wire[15:0] memoryStreamer_io_weights_4;
  wire[15:0] memoryStreamer_io_weights_3;
  wire[15:0] memoryStreamer_io_weights_2;
  wire[15:0] memoryStreamer_io_weights_1;
  wire[15:0] memoryStreamer_io_weights_0;
  wire[7:0] memoryStreamer_io_bias;


  assign T189 = T0[9:0];
  assign T0 = T1;
  assign T1 = {1'h0, Chain_2_io_ys_0};
  assign T190 = T2[9:0];
  assign T2 = T3;
  assign T3 = {1'h0, Chain_2_io_ys_1};
  assign T191 = T4[9:0];
  assign T4 = T5;
  assign T5 = {1'h0, Chain_2_io_ys_2};
  assign T192 = T6[9:0];
  assign T6 = T7;
  assign T7 = {1'h0, Chain_2_io_ys_3};
  assign T193 = T8[9:0];
  assign T8 = T9;
  assign T9 = {1'h0, Chain_2_io_ys_4};
  assign T194 = T10[9:0];
  assign T10 = T11;
  assign T11 = {1'h0, Chain_2_io_ys_5};
  assign T195 = T12[9:0];
  assign T12 = T13;
  assign T13 = {1'h0, Chain_2_io_ys_6};
  assign T196 = T14[9:0];
  assign T14 = T15;
  assign T15 = {1'h0, Chain_2_io_ys_7};
  assign T197 = T16[9:0];
  assign T16 = T17;
  assign T17 = {1'h0, Chain_2_io_ys_8};
  assign T198 = T18[9:0];
  assign T18 = T19;
  assign T19 = {1'h0, Chain_2_io_ys_9};
  assign T199 = T20[9:0];
  assign T20 = T21;
  assign T21 = {1'h0, Chain_2_io_ys_10};
  assign T200 = T22[9:0];
  assign T22 = T23;
  assign T23 = {1'h0, Chain_2_io_ys_11};
  assign T201 = T24[9:0];
  assign T24 = T25;
  assign T25 = {1'h0, Chain_2_io_ys_12};
  assign T202 = T26[9:0];
  assign T26 = T27;
  assign T27 = {1'h0, Chain_2_io_ys_13};
  assign T203 = T28[9:0];
  assign T28 = T29;
  assign T29 = {1'h0, Chain_2_io_ys_14};
  assign T204 = T30[9:0];
  assign T30 = T31;
  assign T31 = {1'h0, Chain_2_io_ys_15};
  assign T205 = T32[9:0];
  assign T32 = T33;
  assign T33 = {1'h0, Chain_1_io_ys_0};
  assign T206 = T34[9:0];
  assign T34 = T35;
  assign T35 = {1'h0, Chain_1_io_ys_1};
  assign T207 = T36[9:0];
  assign T36 = T37;
  assign T37 = {1'h0, Chain_1_io_ys_2};
  assign T208 = T38[9:0];
  assign T38 = T39;
  assign T39 = {1'h0, Chain_1_io_ys_3};
  assign T209 = T40[9:0];
  assign T40 = T41;
  assign T41 = {1'h0, Chain_1_io_ys_4};
  assign T210 = T42[9:0];
  assign T42 = T43;
  assign T43 = {1'h0, Chain_1_io_ys_5};
  assign T211 = T44[9:0];
  assign T44 = T45;
  assign T45 = {1'h0, Chain_1_io_ys_6};
  assign T212 = T46[9:0];
  assign T46 = T47;
  assign T47 = {1'h0, Chain_1_io_ys_7};
  assign T213 = T48[9:0];
  assign T48 = T49;
  assign T49 = {1'h0, Chain_1_io_ys_8};
  assign T214 = T50[9:0];
  assign T50 = T51;
  assign T51 = {1'h0, Chain_1_io_ys_9};
  assign T215 = T52[9:0];
  assign T52 = T53;
  assign T53 = {1'h0, Chain_1_io_ys_10};
  assign T216 = T54[9:0];
  assign T54 = T55;
  assign T55 = {1'h0, Chain_1_io_ys_11};
  assign T217 = T56[9:0];
  assign T56 = T57;
  assign T57 = {1'h0, Chain_1_io_ys_12};
  assign T218 = T58[9:0];
  assign T58 = T59;
  assign T59 = {1'h0, Chain_1_io_ys_13};
  assign T219 = T60[9:0];
  assign T60 = T61;
  assign T61 = {1'h0, Chain_1_io_ys_14};
  assign T220 = T62[9:0];
  assign T62 = T63;
  assign T63 = {1'h0, Chain_1_io_ys_15};
  assign T221 = T64[9:0];
  assign T64 = T65;
  assign T65 = {1'h0, Chain_io_ys_0};
  assign T222 = T66[9:0];
  assign T66 = T67;
  assign T67 = {1'h0, Chain_io_ys_1};
  assign T223 = T68[9:0];
  assign T68 = T69;
  assign T69 = {1'h0, Chain_io_ys_2};
  assign T224 = T70[9:0];
  assign T70 = T71;
  assign T71 = {1'h0, Chain_io_ys_3};
  assign T225 = T72[9:0];
  assign T72 = T73;
  assign T73 = {1'h0, Chain_io_ys_4};
  assign T226 = T74[9:0];
  assign T74 = T75;
  assign T75 = {1'h0, Chain_io_ys_5};
  assign T227 = T76[9:0];
  assign T76 = T77;
  assign T77 = {1'h0, Chain_io_ys_6};
  assign T228 = T78[9:0];
  assign T78 = T79;
  assign T79 = {1'h0, Chain_io_ys_7};
  assign T229 = T80[9:0];
  assign T80 = T81;
  assign T81 = {1'h0, Chain_io_ys_8};
  assign T230 = T82[9:0];
  assign T82 = T83;
  assign T83 = {1'h0, Chain_io_ys_9};
  assign T231 = T84[9:0];
  assign T84 = T85;
  assign T85 = {1'h0, Chain_io_ys_10};
  assign T232 = T86[9:0];
  assign T86 = T87;
  assign T87 = {1'h0, Chain_io_ys_11};
  assign T233 = T88[9:0];
  assign T88 = T89;
  assign T89 = {1'h0, Chain_io_ys_12};
  assign T234 = T90[9:0];
  assign T90 = T91;
  assign T91 = {1'h0, Chain_io_ys_13};
  assign T235 = T92[9:0];
  assign T92 = T93;
  assign T93 = {1'h0, Chain_io_ys_14};
  assign T236 = T94[9:0];
  assign T94 = T95;
  assign T95 = {1'h0, Chain_io_ys_15};
  assign io_done = control_io_done;
  assign io_xOutValid = control_io_valid;
  assign io_xOut_0 = T96;
  assign T96 = T126 ? T112 : T97;
  assign T97 = T111 ? T105 : T98;
  assign T98 = T104 ? T102 : T99;
  assign T99 = T100 ? Activation_io_out_1 : Activation_io_out_0;
  assign T100 = T101[0];
  assign T101 = control_io_selectX;
  assign T102 = T103 ? Activation_io_out_3 : Activation_io_out_2;
  assign T103 = T101[0];
  assign T104 = T101[1];
  assign T105 = T110 ? T108 : T106;
  assign T106 = T107 ? Activation_io_out_5 : Activation_io_out_4;
  assign T107 = T101[0];
  assign T108 = T109 ? Activation_io_out_7 : Activation_io_out_6;
  assign T109 = T101[0];
  assign T110 = T101[1];
  assign T111 = T101[2];
  assign T112 = T125 ? T119 : T113;
  assign T113 = T118 ? T116 : T114;
  assign T114 = T115 ? Activation_io_out_9 : Activation_io_out_8;
  assign T115 = T101[0];
  assign T116 = T117 ? Activation_io_out_11 : Activation_io_out_10;
  assign T117 = T101[0];
  assign T118 = T101[1];
  assign T119 = T124 ? T122 : T120;
  assign T120 = T121 ? Activation_io_out_13 : Activation_io_out_12;
  assign T121 = T101[0];
  assign T122 = T123 ? Activation_io_out_15 : Activation_io_out_14;
  assign T123 = T101[0];
  assign T124 = T101[1];
  assign T125 = T101[2];
  assign T126 = T101[3];
  assign io_xOut_1 = T127;
  assign T127 = T157 ? T143 : T128;
  assign T128 = T142 ? T136 : T129;
  assign T129 = T135 ? T133 : T130;
  assign T130 = T131 ? Activation_1_io_out_1 : Activation_1_io_out_0;
  assign T131 = T132[0];
  assign T132 = control_io_selectX;
  assign T133 = T134 ? Activation_1_io_out_3 : Activation_1_io_out_2;
  assign T134 = T132[0];
  assign T135 = T132[1];
  assign T136 = T141 ? T139 : T137;
  assign T137 = T138 ? Activation_1_io_out_5 : Activation_1_io_out_4;
  assign T138 = T132[0];
  assign T139 = T140 ? Activation_1_io_out_7 : Activation_1_io_out_6;
  assign T140 = T132[0];
  assign T141 = T132[1];
  assign T142 = T132[2];
  assign T143 = T156 ? T150 : T144;
  assign T144 = T149 ? T147 : T145;
  assign T145 = T146 ? Activation_1_io_out_9 : Activation_1_io_out_8;
  assign T146 = T132[0];
  assign T147 = T148 ? Activation_1_io_out_11 : Activation_1_io_out_10;
  assign T148 = T132[0];
  assign T149 = T132[1];
  assign T150 = T155 ? T153 : T151;
  assign T151 = T152 ? Activation_1_io_out_13 : Activation_1_io_out_12;
  assign T152 = T132[0];
  assign T153 = T154 ? Activation_1_io_out_15 : Activation_1_io_out_14;
  assign T154 = T132[0];
  assign T155 = T132[1];
  assign T156 = T132[2];
  assign T157 = T132[3];
  assign io_xOut_2 = T158;
  assign T158 = T188 ? T174 : T159;
  assign T159 = T173 ? T167 : T160;
  assign T160 = T166 ? T164 : T161;
  assign T161 = T162 ? Activation_2_io_out_1 : Activation_2_io_out_0;
  assign T162 = T163[0];
  assign T163 = control_io_selectX;
  assign T164 = T165 ? Activation_2_io_out_3 : Activation_2_io_out_2;
  assign T165 = T163[0];
  assign T166 = T163[1];
  assign T167 = T172 ? T170 : T168;
  assign T168 = T169 ? Activation_2_io_out_5 : Activation_2_io_out_4;
  assign T169 = T163[0];
  assign T170 = T171 ? Activation_2_io_out_7 : Activation_2_io_out_6;
  assign T171 = T163[0];
  assign T172 = T163[1];
  assign T173 = T163[2];
  assign T174 = T187 ? T181 : T175;
  assign T175 = T180 ? T178 : T176;
  assign T176 = T177 ? Activation_2_io_out_9 : Activation_2_io_out_8;
  assign T177 = T163[0];
  assign T178 = T179 ? Activation_2_io_out_11 : Activation_2_io_out_10;
  assign T179 = T163[0];
  assign T180 = T163[1];
  assign T181 = T186 ? T184 : T182;
  assign T182 = T183 ? Activation_2_io_out_13 : Activation_2_io_out_12;
  assign T183 = T163[0];
  assign T184 = T185 ? Activation_2_io_out_15 : Activation_2_io_out_14;
  assign T185 = T163[0];
  assign T186 = T163[1];
  assign T187 = T163[2];
  assign T188 = T163[3];
  assign io_startOut = io_start;
  assign io_ready = control_io_ready;
  WarpControl_1 control(.clk(clk), .reset(reset),
       .io_ready( control_io_ready ),
       .io_start( io_start ),
       .io_nextReady( io_pipeReady ),
       .io_valid( control_io_valid ),
       .io_done( control_io_done ),
       .io_selectX( control_io_selectX ),
       .io_memoryRestart( control_io_memoryRestart ),
       .io_chainRestart( control_io_chainRestart )
  );
  Chain_1 Chain(.clk(clk), .reset(reset),
       .io_weights_15( memoryStreamer_io_weights_15 ),
       .io_weights_14( memoryStreamer_io_weights_14 ),
       .io_weights_13( memoryStreamer_io_weights_13 ),
       .io_weights_12( memoryStreamer_io_weights_12 ),
       .io_weights_11( memoryStreamer_io_weights_11 ),
       .io_weights_10( memoryStreamer_io_weights_10 ),
       .io_weights_9( memoryStreamer_io_weights_9 ),
       .io_weights_8( memoryStreamer_io_weights_8 ),
       .io_weights_7( memoryStreamer_io_weights_7 ),
       .io_weights_6( memoryStreamer_io_weights_6 ),
       .io_weights_5( memoryStreamer_io_weights_5 ),
       .io_weights_4( memoryStreamer_io_weights_4 ),
       .io_weights_3( memoryStreamer_io_weights_3 ),
       .io_weights_2( memoryStreamer_io_weights_2 ),
       .io_weights_1( memoryStreamer_io_weights_1 ),
       .io_weights_0( memoryStreamer_io_weights_0 ),
       .io_bias( memoryStreamer_io_bias ),
       .io_restartIn( control_io_chainRestart ),
       .io_xs( io_xIn_0 ),
       .io_ys_15( Chain_io_ys_15 ),
       .io_ys_14( Chain_io_ys_14 ),
       .io_ys_13( Chain_io_ys_13 ),
       .io_ys_12( Chain_io_ys_12 ),
       .io_ys_11( Chain_io_ys_11 ),
       .io_ys_10( Chain_io_ys_10 ),
       .io_ys_9( Chain_io_ys_9 ),
       .io_ys_8( Chain_io_ys_8 ),
       .io_ys_7( Chain_io_ys_7 ),
       .io_ys_6( Chain_io_ys_6 ),
       .io_ys_5( Chain_io_ys_5 ),
       .io_ys_4( Chain_io_ys_4 ),
       .io_ys_3( Chain_io_ys_3 ),
       .io_ys_2( Chain_io_ys_2 ),
       .io_ys_1( Chain_io_ys_1 ),
       .io_ys_0( Chain_io_ys_0 )
  );
  Chain_1 Chain_1(.clk(clk), .reset(reset),
       .io_weights_15( memoryStreamer_io_weights_15 ),
       .io_weights_14( memoryStreamer_io_weights_14 ),
       .io_weights_13( memoryStreamer_io_weights_13 ),
       .io_weights_12( memoryStreamer_io_weights_12 ),
       .io_weights_11( memoryStreamer_io_weights_11 ),
       .io_weights_10( memoryStreamer_io_weights_10 ),
       .io_weights_9( memoryStreamer_io_weights_9 ),
       .io_weights_8( memoryStreamer_io_weights_8 ),
       .io_weights_7( memoryStreamer_io_weights_7 ),
       .io_weights_6( memoryStreamer_io_weights_6 ),
       .io_weights_5( memoryStreamer_io_weights_5 ),
       .io_weights_4( memoryStreamer_io_weights_4 ),
       .io_weights_3( memoryStreamer_io_weights_3 ),
       .io_weights_2( memoryStreamer_io_weights_2 ),
       .io_weights_1( memoryStreamer_io_weights_1 ),
       .io_weights_0( memoryStreamer_io_weights_0 ),
       .io_bias( memoryStreamer_io_bias ),
       .io_restartIn( control_io_chainRestart ),
       .io_xs( io_xIn_1 ),
       .io_ys_15( Chain_1_io_ys_15 ),
       .io_ys_14( Chain_1_io_ys_14 ),
       .io_ys_13( Chain_1_io_ys_13 ),
       .io_ys_12( Chain_1_io_ys_12 ),
       .io_ys_11( Chain_1_io_ys_11 ),
       .io_ys_10( Chain_1_io_ys_10 ),
       .io_ys_9( Chain_1_io_ys_9 ),
       .io_ys_8( Chain_1_io_ys_8 ),
       .io_ys_7( Chain_1_io_ys_7 ),
       .io_ys_6( Chain_1_io_ys_6 ),
       .io_ys_5( Chain_1_io_ys_5 ),
       .io_ys_4( Chain_1_io_ys_4 ),
       .io_ys_3( Chain_1_io_ys_3 ),
       .io_ys_2( Chain_1_io_ys_2 ),
       .io_ys_1( Chain_1_io_ys_1 ),
       .io_ys_0( Chain_1_io_ys_0 )
  );
  Chain_1 Chain_2(.clk(clk), .reset(reset),
       .io_weights_15( memoryStreamer_io_weights_15 ),
       .io_weights_14( memoryStreamer_io_weights_14 ),
       .io_weights_13( memoryStreamer_io_weights_13 ),
       .io_weights_12( memoryStreamer_io_weights_12 ),
       .io_weights_11( memoryStreamer_io_weights_11 ),
       .io_weights_10( memoryStreamer_io_weights_10 ),
       .io_weights_9( memoryStreamer_io_weights_9 ),
       .io_weights_8( memoryStreamer_io_weights_8 ),
       .io_weights_7( memoryStreamer_io_weights_7 ),
       .io_weights_6( memoryStreamer_io_weights_6 ),
       .io_weights_5( memoryStreamer_io_weights_5 ),
       .io_weights_4( memoryStreamer_io_weights_4 ),
       .io_weights_3( memoryStreamer_io_weights_3 ),
       .io_weights_2( memoryStreamer_io_weights_2 ),
       .io_weights_1( memoryStreamer_io_weights_1 ),
       .io_weights_0( memoryStreamer_io_weights_0 ),
       .io_bias( memoryStreamer_io_bias ),
       .io_restartIn( control_io_chainRestart ),
       .io_xs( io_xIn_2 ),
       .io_ys_15( Chain_2_io_ys_15 ),
       .io_ys_14( Chain_2_io_ys_14 ),
       .io_ys_13( Chain_2_io_ys_13 ),
       .io_ys_12( Chain_2_io_ys_12 ),
       .io_ys_11( Chain_2_io_ys_11 ),
       .io_ys_10( Chain_2_io_ys_10 ),
       .io_ys_9( Chain_2_io_ys_9 ),
       .io_ys_8( Chain_2_io_ys_8 ),
       .io_ys_7( Chain_2_io_ys_7 ),
       .io_ys_6( Chain_2_io_ys_6 ),
       .io_ys_5( Chain_2_io_ys_5 ),
       .io_ys_4( Chain_2_io_ys_4 ),
       .io_ys_3( Chain_2_io_ys_3 ),
       .io_ys_2( Chain_2_io_ys_2 ),
       .io_ys_1( Chain_2_io_ys_1 ),
       .io_ys_0( Chain_2_io_ys_0 )
  );
  Activation_1 Activation(
       .io_in_15( T236 ),
       .io_in_14( T235 ),
       .io_in_13( T234 ),
       .io_in_12( T233 ),
       .io_in_11( T232 ),
       .io_in_10( T231 ),
       .io_in_9( T230 ),
       .io_in_8( T229 ),
       .io_in_7( T228 ),
       .io_in_6( T227 ),
       .io_in_5( T226 ),
       .io_in_4( T225 ),
       .io_in_3( T224 ),
       .io_in_2( T223 ),
       .io_in_1( T222 ),
       .io_in_0( T221 ),
       .io_out_15( Activation_io_out_15 ),
       .io_out_14( Activation_io_out_14 ),
       .io_out_13( Activation_io_out_13 ),
       .io_out_12( Activation_io_out_12 ),
       .io_out_11( Activation_io_out_11 ),
       .io_out_10( Activation_io_out_10 ),
       .io_out_9( Activation_io_out_9 ),
       .io_out_8( Activation_io_out_8 ),
       .io_out_7( Activation_io_out_7 ),
       .io_out_6( Activation_io_out_6 ),
       .io_out_5( Activation_io_out_5 ),
       .io_out_4( Activation_io_out_4 ),
       .io_out_3( Activation_io_out_3 ),
       .io_out_2( Activation_io_out_2 ),
       .io_out_1( Activation_io_out_1 ),
       .io_out_0( Activation_io_out_0 )
  );
  Activation_1 Activation_1(
       .io_in_15( T220 ),
       .io_in_14( T219 ),
       .io_in_13( T218 ),
       .io_in_12( T217 ),
       .io_in_11( T216 ),
       .io_in_10( T215 ),
       .io_in_9( T214 ),
       .io_in_8( T213 ),
       .io_in_7( T212 ),
       .io_in_6( T211 ),
       .io_in_5( T210 ),
       .io_in_4( T209 ),
       .io_in_3( T208 ),
       .io_in_2( T207 ),
       .io_in_1( T206 ),
       .io_in_0( T205 ),
       .io_out_15( Activation_1_io_out_15 ),
       .io_out_14( Activation_1_io_out_14 ),
       .io_out_13( Activation_1_io_out_13 ),
       .io_out_12( Activation_1_io_out_12 ),
       .io_out_11( Activation_1_io_out_11 ),
       .io_out_10( Activation_1_io_out_10 ),
       .io_out_9( Activation_1_io_out_9 ),
       .io_out_8( Activation_1_io_out_8 ),
       .io_out_7( Activation_1_io_out_7 ),
       .io_out_6( Activation_1_io_out_6 ),
       .io_out_5( Activation_1_io_out_5 ),
       .io_out_4( Activation_1_io_out_4 ),
       .io_out_3( Activation_1_io_out_3 ),
       .io_out_2( Activation_1_io_out_2 ),
       .io_out_1( Activation_1_io_out_1 ),
       .io_out_0( Activation_1_io_out_0 )
  );
  Activation_1 Activation_2(
       .io_in_15( T204 ),
       .io_in_14( T203 ),
       .io_in_13( T202 ),
       .io_in_12( T201 ),
       .io_in_11( T200 ),
       .io_in_10( T199 ),
       .io_in_9( T198 ),
       .io_in_8( T197 ),
       .io_in_7( T196 ),
       .io_in_6( T195 ),
       .io_in_5( T194 ),
       .io_in_4( T193 ),
       .io_in_3( T192 ),
       .io_in_2( T191 ),
       .io_in_1( T190 ),
       .io_in_0( T189 ),
       .io_out_15( Activation_2_io_out_15 ),
       .io_out_14( Activation_2_io_out_14 ),
       .io_out_13( Activation_2_io_out_13 ),
       .io_out_12( Activation_2_io_out_12 ),
       .io_out_11( Activation_2_io_out_11 ),
       .io_out_10( Activation_2_io_out_10 ),
       .io_out_9( Activation_2_io_out_9 ),
       .io_out_8( Activation_2_io_out_8 ),
       .io_out_7( Activation_2_io_out_7 ),
       .io_out_6( Activation_2_io_out_6 ),
       .io_out_5( Activation_2_io_out_5 ),
       .io_out_4( Activation_2_io_out_4 ),
       .io_out_3( Activation_2_io_out_3 ),
       .io_out_2( Activation_2_io_out_2 ),
       .io_out_1( Activation_2_io_out_1 ),
       .io_out_0( Activation_2_io_out_0 )
  );
  MemoryStreamer_2 memoryStreamer(.clk(clk), .reset(reset),
       .io_restart( control_io_memoryRestart ),
       .io_weights_15( memoryStreamer_io_weights_15 ),
       .io_weights_14( memoryStreamer_io_weights_14 ),
       .io_weights_13( memoryStreamer_io_weights_13 ),
       .io_weights_12( memoryStreamer_io_weights_12 ),
       .io_weights_11( memoryStreamer_io_weights_11 ),
       .io_weights_10( memoryStreamer_io_weights_10 ),
       .io_weights_9( memoryStreamer_io_weights_9 ),
       .io_weights_8( memoryStreamer_io_weights_8 ),
       .io_weights_7( memoryStreamer_io_weights_7 ),
       .io_weights_6( memoryStreamer_io_weights_6 ),
       .io_weights_5( memoryStreamer_io_weights_5 ),
       .io_weights_4( memoryStreamer_io_weights_4 ),
       .io_weights_3( memoryStreamer_io_weights_3 ),
       .io_weights_2( memoryStreamer_io_weights_2 ),
       .io_weights_1( memoryStreamer_io_weights_1 ),
       .io_weights_0( memoryStreamer_io_weights_0 ),
       .io_bias( memoryStreamer_io_bias )
  );
endmodule

module WarpControl_2(input clk, input reset,
    output io_ready,
    input  io_start,
    input  io_nextReady,
    output io_valid,
    output io_done,
    output[3:0] io_selectX,
    output io_memoryRestart,
    output io_chainRestart
);

  wire signalDone;
  reg  signalTailing;
  wire T8;
  wire signalLastActiveCycle;
  wire signalResetSelectX;
  reg  signalFirstOutputCycle;
  wire T9;
  wire signalOutputtingNext;
  wire T0;
  wire signalFirstReadyCycle;
  wire T1;
  wire signalLastCycleInPass;
  wire signalStartNewPass;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire[3:0] cycleInPass_io_value;
  wire[3:0] cycle_io_value;
  wire[3:0] tailCycle_io_value;
  wire[3:0] selectX_io_value;
  wire isActive_io_state;
  wire isReady_io_state;
  wire isOutputting_io_state;
  wire isTailing_io_state;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    signalTailing = {1{$random}};
    signalFirstOutputCycle = {1{$random}};
  end
// synthesis translate_on
`endif

  assign signalDone = tailCycle_io_value == 4'h9;
  assign T8 = reset ? 1'h0 : signalLastActiveCycle;
  assign signalLastActiveCycle = cycle_io_value == 4'hf;
  assign signalResetSelectX = selectX_io_value == 4'h9;
  assign T9 = reset ? 1'h0 : signalOutputtingNext;
  assign signalOutputtingNext = T0 & isActive_io_state;
  assign T0 = cycleInPass_io_value == 4'hf;
  assign signalFirstReadyCycle = T1 & isTailing_io_state;
  assign T1 = tailCycle_io_value == 4'h0;
  assign signalLastCycleInPass = cycleInPass_io_value == 4'hf;
  assign io_chainRestart = signalStartNewPass;
  assign signalStartNewPass = cycleInPass_io_value == 4'h0;
  assign io_memoryRestart = T2;
  assign T2 = T4 & T3;
  assign T3 = io_start ^ 1'h1;
  assign T4 = isReady_io_state | signalLastActiveCycle;
  assign io_selectX = selectX_io_value;
  assign io_done = signalDone;
  assign io_valid = isOutputting_io_state;
  assign io_ready = T5;
  assign T5 = T7 & T6;
  assign T6 = io_start ^ 1'h1;
  assign T7 = isReady_io_state & io_nextReady;
  Counter_2 cycleInPass(.clk(clk), .reset(reset),
       .io_enable( isActive_io_state ),
       .io_rst( signalLastCycleInPass ),
       .io_value( cycleInPass_io_value )
  );
  Counter_2 cycle(.clk(clk), .reset(reset),
       .io_enable( isActive_io_state ),
       .io_rst( signalLastActiveCycle ),
       .io_value( cycle_io_value )
  );
  Counter_2 tailCycle(.clk(clk), .reset(reset),
       .io_enable( isTailing_io_state ),
       .io_rst( signalDone ),
       .io_value( tailCycle_io_value )
  );
  Counter_2 selectX(.clk(clk), .reset(reset),
       .io_enable( isOutputting_io_state ),
       .io_rst( signalResetSelectX ),
       .io_value( selectX_io_value )
  );
  Switch_0 isActive(.clk(clk), .reset(reset),
       .io_signalOn( io_start ),
       .io_state( isActive_io_state ),
       .io_rst( signalLastActiveCycle )
  );
  Switch_1 isReady(.clk(clk), .reset(reset),
       .io_signalOn( signalFirstReadyCycle ),
       .io_state( isReady_io_state ),
       .io_rst( io_start )
  );
  Switch_0 isOutputting(.clk(clk), .reset(reset),
       .io_signalOn( signalFirstOutputCycle ),
       .io_state( isOutputting_io_state ),
       .io_rst( signalResetSelectX )
  );
  Switch_0 isTailing(.clk(clk), .reset(reset),
       .io_signalOn( signalTailing ),
       .io_state( isTailing_io_state ),
       .io_rst( signalDone )
  );

  always @(posedge clk) begin
    if(reset) begin
      signalTailing <= 1'h0;
    end else begin
      signalTailing <= signalLastActiveCycle;
    end
    if(reset) begin
      signalFirstOutputCycle <= 1'h0;
    end else begin
      signalFirstOutputCycle <= signalOutputtingNext;
    end
  end
endmodule

module Chain_2(input clk, input reset,
    input [15:0] io_weights_9,
    input [15:0] io_weights_8,
    input [15:0] io_weights_7,
    input [15:0] io_weights_6,
    input [15:0] io_weights_5,
    input [15:0] io_weights_4,
    input [15:0] io_weights_3,
    input [15:0] io_weights_2,
    input [15:0] io_weights_1,
    input [15:0] io_weights_0,
    input [7:0] io_bias,
    input  io_restartIn,
    input [15:0] io_xs,
    output[9:0] io_ys_9,
    output[9:0] io_ys_8,
    output[9:0] io_ys_7,
    output[9:0] io_ys_6,
    output[9:0] io_ys_5,
    output[9:0] io_ys_4,
    output[9:0] io_ys_3,
    output[9:0] io_ys_2,
    output[9:0] io_ys_1,
    output[9:0] io_ys_0
);

  wire[7:0] T20;
  wire[8:0] T0;
  wire[8:0] T1;
  wire[7:0] T21;
  wire[8:0] T2;
  wire[8:0] T3;
  wire[7:0] T22;
  wire[8:0] T4;
  wire[8:0] T5;
  wire[7:0] T23;
  wire[8:0] T6;
  wire[8:0] T7;
  wire[7:0] T24;
  wire[8:0] T8;
  wire[8:0] T9;
  wire[7:0] T25;
  wire[8:0] T10;
  wire[8:0] T11;
  wire[7:0] T26;
  wire[8:0] T12;
  wire[8:0] T13;
  wire[7:0] T27;
  wire[8:0] T14;
  wire[8:0] T15;
  wire[7:0] T28;
  wire[8:0] T16;
  wire[8:0] T17;
  wire[7:0] T29;
  wire[8:0] T18;
  wire[8:0] T19;
  wire[15:0] ProcessingUnit_io_xOut;
  wire[9:0] ProcessingUnit_io_yOut;
  wire ProcessingUnit_io_restartOut;
  wire[15:0] ProcessingUnit_1_io_xOut;
  wire[9:0] ProcessingUnit_1_io_yOut;
  wire ProcessingUnit_1_io_restartOut;
  wire[15:0] ProcessingUnit_2_io_xOut;
  wire[9:0] ProcessingUnit_2_io_yOut;
  wire ProcessingUnit_2_io_restartOut;
  wire[15:0] ProcessingUnit_3_io_xOut;
  wire[9:0] ProcessingUnit_3_io_yOut;
  wire ProcessingUnit_3_io_restartOut;
  wire[15:0] ProcessingUnit_4_io_xOut;
  wire[9:0] ProcessingUnit_4_io_yOut;
  wire ProcessingUnit_4_io_restartOut;
  wire[15:0] ProcessingUnit_5_io_xOut;
  wire[9:0] ProcessingUnit_5_io_yOut;
  wire ProcessingUnit_5_io_restartOut;
  wire[15:0] ProcessingUnit_6_io_xOut;
  wire[9:0] ProcessingUnit_6_io_yOut;
  wire ProcessingUnit_6_io_restartOut;
  wire[15:0] ProcessingUnit_7_io_xOut;
  wire[9:0] ProcessingUnit_7_io_yOut;
  wire ProcessingUnit_7_io_restartOut;
  wire[15:0] ProcessingUnit_8_io_xOut;
  wire[9:0] ProcessingUnit_8_io_yOut;
  wire ProcessingUnit_8_io_restartOut;
  wire[9:0] ProcessingUnit_9_io_yOut;


  assign T20 = T0[7:0];
  assign T0 = T1;
  assign T1 = {1'h0, io_bias};
  assign T21 = T2[7:0];
  assign T2 = T3;
  assign T3 = {1'h0, io_bias};
  assign T22 = T4[7:0];
  assign T4 = T5;
  assign T5 = {1'h0, io_bias};
  assign T23 = T6[7:0];
  assign T6 = T7;
  assign T7 = {1'h0, io_bias};
  assign T24 = T8[7:0];
  assign T8 = T9;
  assign T9 = {1'h0, io_bias};
  assign T25 = T10[7:0];
  assign T10 = T11;
  assign T11 = {1'h0, io_bias};
  assign T26 = T12[7:0];
  assign T12 = T13;
  assign T13 = {1'h0, io_bias};
  assign T27 = T14[7:0];
  assign T14 = T15;
  assign T15 = {1'h0, io_bias};
  assign T28 = T16[7:0];
  assign T16 = T17;
  assign T17 = {1'h0, io_bias};
  assign T29 = T18[7:0];
  assign T18 = T19;
  assign T19 = {1'h0, io_bias};
  assign io_ys_0 = ProcessingUnit_io_yOut;
  assign io_ys_1 = ProcessingUnit_1_io_yOut;
  assign io_ys_2 = ProcessingUnit_2_io_yOut;
  assign io_ys_3 = ProcessingUnit_3_io_yOut;
  assign io_ys_4 = ProcessingUnit_4_io_yOut;
  assign io_ys_5 = ProcessingUnit_5_io_yOut;
  assign io_ys_6 = ProcessingUnit_6_io_yOut;
  assign io_ys_7 = ProcessingUnit_7_io_yOut;
  assign io_ys_8 = ProcessingUnit_8_io_yOut;
  assign io_ys_9 = ProcessingUnit_9_io_yOut;
  ProcessingUnit ProcessingUnit(.clk(clk), .reset(reset),
       .io_xs( io_xs ),
       .io_ws( io_weights_0 ),
       .io_xOut( ProcessingUnit_io_xOut ),
       .io_yOut( ProcessingUnit_io_yOut ),
       .io_bias( T29 ),
       .io_restartIn( io_restartIn ),
       .io_restartOut( ProcessingUnit_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_1(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_io_xOut ),
       .io_ws( io_weights_1 ),
       .io_xOut( ProcessingUnit_1_io_xOut ),
       .io_yOut( ProcessingUnit_1_io_yOut ),
       .io_bias( T28 ),
       .io_restartIn( ProcessingUnit_io_restartOut ),
       .io_restartOut( ProcessingUnit_1_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_2(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_1_io_xOut ),
       .io_ws( io_weights_2 ),
       .io_xOut( ProcessingUnit_2_io_xOut ),
       .io_yOut( ProcessingUnit_2_io_yOut ),
       .io_bias( T27 ),
       .io_restartIn( ProcessingUnit_1_io_restartOut ),
       .io_restartOut( ProcessingUnit_2_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_3(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_2_io_xOut ),
       .io_ws( io_weights_3 ),
       .io_xOut( ProcessingUnit_3_io_xOut ),
       .io_yOut( ProcessingUnit_3_io_yOut ),
       .io_bias( T26 ),
       .io_restartIn( ProcessingUnit_2_io_restartOut ),
       .io_restartOut( ProcessingUnit_3_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_4(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_3_io_xOut ),
       .io_ws( io_weights_4 ),
       .io_xOut( ProcessingUnit_4_io_xOut ),
       .io_yOut( ProcessingUnit_4_io_yOut ),
       .io_bias( T25 ),
       .io_restartIn( ProcessingUnit_3_io_restartOut ),
       .io_restartOut( ProcessingUnit_4_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_5(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_4_io_xOut ),
       .io_ws( io_weights_5 ),
       .io_xOut( ProcessingUnit_5_io_xOut ),
       .io_yOut( ProcessingUnit_5_io_yOut ),
       .io_bias( T24 ),
       .io_restartIn( ProcessingUnit_4_io_restartOut ),
       .io_restartOut( ProcessingUnit_5_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_6(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_5_io_xOut ),
       .io_ws( io_weights_6 ),
       .io_xOut( ProcessingUnit_6_io_xOut ),
       .io_yOut( ProcessingUnit_6_io_yOut ),
       .io_bias( T23 ),
       .io_restartIn( ProcessingUnit_5_io_restartOut ),
       .io_restartOut( ProcessingUnit_6_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_7(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_6_io_xOut ),
       .io_ws( io_weights_7 ),
       .io_xOut( ProcessingUnit_7_io_xOut ),
       .io_yOut( ProcessingUnit_7_io_yOut ),
       .io_bias( T22 ),
       .io_restartIn( ProcessingUnit_6_io_restartOut ),
       .io_restartOut( ProcessingUnit_7_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_8(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_7_io_xOut ),
       .io_ws( io_weights_8 ),
       .io_xOut( ProcessingUnit_8_io_xOut ),
       .io_yOut( ProcessingUnit_8_io_yOut ),
       .io_bias( T21 ),
       .io_restartIn( ProcessingUnit_7_io_restartOut ),
       .io_restartOut( ProcessingUnit_8_io_restartOut )
  );
  ProcessingUnit ProcessingUnit_9(.clk(clk), .reset(reset),
       .io_xs( ProcessingUnit_8_io_xOut ),
       .io_ws( io_weights_9 ),
       //.io_xOut(  )
       .io_yOut( ProcessingUnit_9_io_yOut ),
       .io_bias( T20 ),
       .io_restartIn( ProcessingUnit_8_io_restartOut )
       //.io_restartOut(  )
  );
endmodule

module Activation_2(
    input [9:0] io_in_9,
    input [9:0] io_in_8,
    input [9:0] io_in_7,
    input [9:0] io_in_6,
    input [9:0] io_in_5,
    input [9:0] io_in_4,
    input [9:0] io_in_3,
    input [9:0] io_in_2,
    input [9:0] io_in_1,
    input [9:0] io_in_0,
    output io_out_9,
    output io_out_8,
    output io_out_7,
    output io_out_6,
    output io_out_5,
    output io_out_4,
    output io_out_3,
    output io_out_2,
    output io_out_1,
    output io_out_0
);

  wire T0;
  wire T1;
  wire[12:0] T2;
  wire[12:0] T3;
  wire T4;
  wire T5;
  wire[12:0] T6;
  wire[12:0] T7;
  wire T8;
  wire T9;
  wire[12:0] T10;
  wire[12:0] T11;
  wire T12;
  wire T13;
  wire[12:0] T14;
  wire[12:0] T15;
  wire T16;
  wire T17;
  wire[12:0] T18;
  wire[12:0] T19;
  wire T20;
  wire T21;
  wire[12:0] T22;
  wire[12:0] T23;
  wire T24;
  wire T25;
  wire[12:0] T26;
  wire[12:0] T27;
  wire T28;
  wire T29;
  wire[12:0] T30;
  wire[12:0] T31;
  wire T32;
  wire T33;
  wire[12:0] T34;
  wire[12:0] T35;
  wire T36;
  wire T37;
  wire[12:0] T38;
  wire[12:0] T39;


  assign io_out_0 = T0;
  assign T0 = ~ T1;
  assign T1 = T2[9];
  assign T2 = T3 - 13'h100;
  assign T3 = $signed(io_in_0) * $signed(3'h2);
  assign io_out_1 = T4;
  assign T4 = ~ T5;
  assign T5 = T6[9];
  assign T6 = T7 - 13'h100;
  assign T7 = $signed(io_in_1) * $signed(3'h2);
  assign io_out_2 = T8;
  assign T8 = ~ T9;
  assign T9 = T10[9];
  assign T10 = T11 - 13'h100;
  assign T11 = $signed(io_in_2) * $signed(3'h2);
  assign io_out_3 = T12;
  assign T12 = ~ T13;
  assign T13 = T14[9];
  assign T14 = T15 - 13'h100;
  assign T15 = $signed(io_in_3) * $signed(3'h2);
  assign io_out_4 = T16;
  assign T16 = ~ T17;
  assign T17 = T18[9];
  assign T18 = T19 - 13'h100;
  assign T19 = $signed(io_in_4) * $signed(3'h2);
  assign io_out_5 = T20;
  assign T20 = ~ T21;
  assign T21 = T22[9];
  assign T22 = T23 - 13'h100;
  assign T23 = $signed(io_in_5) * $signed(3'h2);
  assign io_out_6 = T24;
  assign T24 = ~ T25;
  assign T25 = T26[9];
  assign T26 = T27 - 13'h100;
  assign T27 = $signed(io_in_6) * $signed(3'h2);
  assign io_out_7 = T28;
  assign T28 = ~ T29;
  assign T29 = T30[9];
  assign T30 = T31 - 13'h100;
  assign T31 = $signed(io_in_7) * $signed(3'h2);
  assign io_out_8 = T32;
  assign T32 = ~ T33;
  assign T33 = T34[9];
  assign T34 = T35 - 13'h100;
  assign T35 = $signed(io_in_8) * $signed(3'h2);
  assign io_out_9 = T36;
  assign T36 = ~ T37;
  assign T37 = T38[9];
  assign T38 = T39 - 13'h100;
  assign T39 = $signed(io_in_9) * $signed(3'h2);
endmodule

module MemoryUnit_35(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[3:0] T5;
  wire[4:0] addr;
  reg [4:0] counter;
  wire[4:0] T6;
  wire[4:0] T2;
  wire[4:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (T5)
    0: T0 = 32'hc24f5e78;
    1: T0 = 32'h35871eb5;
    2: T0 = 32'hf043786a;
    3: T0 = 32'hc701ec94;
    4: T0 = 32'h1221d7da;
    5: T0 = 32'hb30548e8;
    6: T0 = 32'h3b1ba226;
    7: T0 = 32'h7478163d;
    8: T0 = 32'h8bc67614;
    9: T0 = 32'he9fd3d40;
    10: T0 = 32'h47be126e;
    11: T0 = 32'hefb3058a;
    12: T0 = 32'h3f65c8a1;
    13: T0 = 32'ha766e982;
    14: T0 = 32'h9658a1bf;
    15: T0 = 32'h16493133;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[3:0];
  assign addr = io_restartIn ? 5'h0 : counter;
  assign T6 = reset ? 5'h0 : T2;
  assign T2 = io_restartIn ? 5'h1 : T3;
  assign T3 = counter + 5'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 5'h0;
    end else if(io_restartIn) begin
      counter <= 5'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_36(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[3:0] T5;
  wire[4:0] addr;
  reg [4:0] counter;
  wire[4:0] T6;
  wire[4:0] T2;
  wire[4:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (T5)
    0: T0 = 32'hce327169;
    1: T0 = 32'haca6720e;
    2: T0 = 32'h8c1a3cd8;
    3: T0 = 32'h3acf6236;
    4: T0 = 32'h21bd644b;
    5: T0 = 32'hf9c77753;
    6: T0 = 32'ha44d8ecd;
    7: T0 = 32'h5108944f;
    8: T0 = 32'h6a0cf020;
    9: T0 = 32'he31ea5ab;
    10: T0 = 32'hda031a1e;
    11: T0 = 32'h4575d931;
    12: T0 = 32'h88fea3da;
    13: T0 = 32'hf345197d;
    14: T0 = 32'he3ecbba5;
    15: T0 = 32'he6705606;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[3:0];
  assign addr = io_restartIn ? 5'h0 : counter;
  assign T6 = reset ? 5'h0 : T2;
  assign T2 = io_restartIn ? 5'h1 : T3;
  assign T3 = counter + 5'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 5'h0;
    end else if(io_restartIn) begin
      counter <= 5'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_37(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[3:0] T5;
  wire[4:0] addr;
  reg [4:0] counter;
  wire[4:0] T6;
  wire[4:0] T2;
  wire[4:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (T5)
    0: T0 = 32'hc1f1261e;
    1: T0 = 32'he3f4fe62;
    2: T0 = 32'hdb1fadb7;
    3: T0 = 32'he0c7eac6;
    4: T0 = 32'hbaf1173a;
    5: T0 = 32'ha46cddf7;
    6: T0 = 32'h82a4d217;
    7: T0 = 32'h8993f837;
    8: T0 = 32'h65ec5eb2;
    9: T0 = 32'h88d4fddb;
    10: T0 = 32'hcab6b913;
    11: T0 = 32'ha7e43a78;
    12: T0 = 32'ha195ac16;
    13: T0 = 32'h4ec78676;
    14: T0 = 32'h23abf796;
    15: T0 = 32'h882e2cdf;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[3:0];
  assign addr = io_restartIn ? 5'h0 : counter;
  assign T6 = reset ? 5'h0 : T2;
  assign T2 = io_restartIn ? 5'h1 : T3;
  assign T3 = counter + 5'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 5'h0;
    end else if(io_restartIn) begin
      counter <= 5'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_38(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[3:0] T5;
  wire[4:0] addr;
  reg [4:0] counter;
  wire[4:0] T6;
  wire[4:0] T2;
  wire[4:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (T5)
    0: T0 = 32'hb52cc899;
    1: T0 = 32'hde69bdb1;
    2: T0 = 32'hb46c020;
    3: T0 = 32'h9f6d956a;
    4: T0 = 32'h694f0031;
    5: T0 = 32'ha9d556ee;
    6: T0 = 32'hbb128f17;
    7: T0 = 32'h63e19481;
    8: T0 = 32'h29722489;
    9: T0 = 32'h177f4524;
    10: T0 = 32'hb2d6be4d;
    11: T0 = 32'h4992aed6;
    12: T0 = 32'hc36917af;
    13: T0 = 32'h44109f87;
    14: T0 = 32'h78390b81;
    15: T0 = 32'h75ff28c4;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[3:0];
  assign addr = io_restartIn ? 5'h0 : counter;
  assign T6 = reset ? 5'h0 : T2;
  assign T2 = io_restartIn ? 5'h1 : T3;
  assign T3 = counter + 5'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 5'h0;
    end else if(io_restartIn) begin
      counter <= 5'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_39(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[31:0] io_weights
);

  reg [31:0] weightsReg;
  wire[31:0] T4;
  reg [31:0] T0;
  wire[3:0] T5;
  wire[4:0] addr;
  reg [4:0] counter;
  wire[4:0] T6;
  wire[4:0] T2;
  wire[4:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 32'h0 : T0;
  always @(*) case (T5)
    0: T0 = 32'h2adb055c;
    1: T0 = 32'h8b8704ed;
    2: T0 = 32'hc179e371;
    3: T0 = 32'h1f96d38e;
    4: T0 = 32'h1cc98c2d;
    5: T0 = 32'h1cf02ccb;
    6: T0 = 32'hcc24b4d8;
    7: T0 = 32'h5ce876f1;
    8: T0 = 32'hf50aafab;
    9: T0 = 32'h5b63cc27;
    10: T0 = 32'h325930ec;
    11: T0 = 32'he5f950ab;
    12: T0 = 32'h768e18f0;
    13: T0 = 32'h59b9449f;
    14: T0 = 32'hfc803110;
    15: T0 = 32'h4c8a7fbd;
    default: begin
      T0 = 32'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[3:0];
  assign addr = io_restartIn ? 5'h0 : counter;
  assign T6 = reset ? 5'h0 : T2;
  assign T2 = io_restartIn ? 5'h1 : T3;
  assign T3 = counter + 5'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 32'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 5'h0;
    end else if(io_restartIn) begin
      counter <= 5'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryUnit_40(input clk, input reset,
    input  io_restartIn,
    output io_restartOut,
    output[7:0] io_weights
);

  reg [7:0] weightsReg;
  wire[7:0] T4;
  reg [7:0] T0;
  wire[3:0] T5;
  wire[4:0] addr;
  reg [4:0] counter;
  wire[4:0] T6;
  wire[4:0] T2;
  wire[4:0] T3;
  reg  restartRegs_1;
  wire T7;
  reg  restartRegs_0;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    weightsReg = {1{$random}};
    counter = {1{$random}};
    restartRegs_1 = {1{$random}};
    restartRegs_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_weights = weightsReg;
  assign T4 = reset ? 8'h0 : T0;
  always @(*) case (T5)
    0: T0 = 8'hc6;
    1: T0 = 8'hc9;
    2: T0 = 8'hc5;
    3: T0 = 8'hc9;
    4: T0 = 8'hca;
    5: T0 = 8'hc9;
    6: T0 = 8'hc7;
    7: T0 = 8'hcb;
    8: T0 = 8'hc9;
    9: T0 = 8'hc8;
    10: T0 = 8'h0;
    11: T0 = 8'h0;
    12: T0 = 8'h0;
    13: T0 = 8'h0;
    14: T0 = 8'h0;
    15: T0 = 8'h0;
    default: begin
      T0 = 8'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T0 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T5 = addr[3:0];
  assign addr = io_restartIn ? 5'h0 : counter;
  assign T6 = reset ? 5'h0 : T2;
  assign T2 = io_restartIn ? 5'h1 : T3;
  assign T3 = counter + 5'h1;
  assign io_restartOut = restartRegs_1;
  assign T7 = reset ? 1'h0 : restartRegs_0;
  assign T8 = reset ? 1'h0 : io_restartIn;

  always @(posedge clk) begin
    if(reset) begin
      weightsReg <= 8'h0;
    end else begin
      weightsReg <= T0;
    end
    if(reset) begin
      counter <= 5'h0;
    end else if(io_restartIn) begin
      counter <= 5'h1;
    end else begin
      counter <= T3;
    end
    if(reset) begin
      restartRegs_1 <= 1'h0;
    end else begin
      restartRegs_1 <= restartRegs_0;
    end
    if(reset) begin
      restartRegs_0 <= 1'h0;
    end else begin
      restartRegs_0 <= io_restartIn;
    end
  end
endmodule

module MemoryStreamer_3(input clk, input reset,
    input  io_restart,
    output[15:0] io_weights_9,
    output[15:0] io_weights_8,
    output[15:0] io_weights_7,
    output[15:0] io_weights_6,
    output[15:0] io_weights_5,
    output[15:0] io_weights_4,
    output[15:0] io_weights_3,
    output[15:0] io_weights_2,
    output[15:0] io_weights_1,
    output[15:0] io_weights_0,
    output[7:0] io_bias
);

  wire[7:0] T12;
  wire[8:0] T0;
  wire[8:0] T1;
  wire[15:0] T2;
  wire[15:0] T3;
  wire[15:0] T4;
  wire[15:0] T5;
  wire[15:0] T6;
  wire[15:0] T7;
  wire[15:0] T8;
  wire[15:0] T9;
  wire[15:0] T10;
  wire[15:0] T11;
  wire MemoryUnit_io_restartOut;
  wire[31:0] MemoryUnit_io_weights;
  wire MemoryUnit_1_io_restartOut;
  wire[31:0] MemoryUnit_1_io_weights;
  wire MemoryUnit_2_io_restartOut;
  wire[31:0] MemoryUnit_2_io_weights;
  wire MemoryUnit_3_io_restartOut;
  wire[31:0] MemoryUnit_3_io_weights;
  wire[31:0] MemoryUnit_4_io_weights;
  wire[7:0] biasMemoryUnit_io_weights;


  assign io_bias = T12;
  assign T12 = T0[7:0];
  assign T0 = T1;
  assign T1 = {1'h0, biasMemoryUnit_io_weights};
  assign io_weights_0 = T2;
  assign T2 = MemoryUnit_io_weights[15:0];
  assign io_weights_1 = T3;
  assign T3 = MemoryUnit_io_weights[31:16];
  assign io_weights_2 = T4;
  assign T4 = MemoryUnit_1_io_weights[15:0];
  assign io_weights_3 = T5;
  assign T5 = MemoryUnit_1_io_weights[31:16];
  assign io_weights_4 = T6;
  assign T6 = MemoryUnit_2_io_weights[15:0];
  assign io_weights_5 = T7;
  assign T7 = MemoryUnit_2_io_weights[31:16];
  assign io_weights_6 = T8;
  assign T8 = MemoryUnit_3_io_weights[15:0];
  assign io_weights_7 = T9;
  assign T9 = MemoryUnit_3_io_weights[31:16];
  assign io_weights_8 = T10;
  assign T10 = MemoryUnit_4_io_weights[15:0];
  assign io_weights_9 = T11;
  assign T11 = MemoryUnit_4_io_weights[31:16];
  MemoryUnit_35 MemoryUnit(.clk(clk), .reset(reset),
       .io_restartIn( io_restart ),
       .io_restartOut( MemoryUnit_io_restartOut ),
       .io_weights( MemoryUnit_io_weights )
  );
  MemoryUnit_36 MemoryUnit_1(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_io_restartOut ),
       .io_restartOut( MemoryUnit_1_io_restartOut ),
       .io_weights( MemoryUnit_1_io_weights )
  );
  MemoryUnit_37 MemoryUnit_2(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_1_io_restartOut ),
       .io_restartOut( MemoryUnit_2_io_restartOut ),
       .io_weights( MemoryUnit_2_io_weights )
  );
  MemoryUnit_38 MemoryUnit_3(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_2_io_restartOut ),
       .io_restartOut( MemoryUnit_3_io_restartOut ),
       .io_weights( MemoryUnit_3_io_weights )
  );
  MemoryUnit_39 MemoryUnit_4(.clk(clk), .reset(reset),
       .io_restartIn( MemoryUnit_3_io_restartOut ),
       //.io_restartOut(  )
       .io_weights( MemoryUnit_4_io_weights )
  );
  MemoryUnit_40 biasMemoryUnit(.clk(clk), .reset(reset),
       .io_restartIn( io_restart ),
       //.io_restartOut(  )
       .io_weights( biasMemoryUnit_io_weights )
  );
endmodule

module Warp_3(input clk, input reset,
    input [15:0] io_xIn_0,
    input  io_start,
    output io_ready,
    output io_startOut,
    output io_xOut_0,
    output io_xOutValid,
    input  io_pipeReady,
    output io_done
);

  wire[9:0] T39;
  wire[10:0] T0;
  wire[10:0] T1;
  wire[9:0] T40;
  wire[10:0] T2;
  wire[10:0] T3;
  wire[9:0] T41;
  wire[10:0] T4;
  wire[10:0] T5;
  wire[9:0] T42;
  wire[10:0] T6;
  wire[10:0] T7;
  wire[9:0] T43;
  wire[10:0] T8;
  wire[10:0] T9;
  wire[9:0] T44;
  wire[10:0] T10;
  wire[10:0] T11;
  wire[9:0] T45;
  wire[10:0] T12;
  wire[10:0] T13;
  wire[9:0] T46;
  wire[10:0] T14;
  wire[10:0] T15;
  wire[9:0] T47;
  wire[10:0] T16;
  wire[10:0] T17;
  wire[9:0] T48;
  wire[10:0] T18;
  wire[10:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[3:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire Activation_io_out_9;
  wire Activation_io_out_8;
  wire Activation_io_out_7;
  wire Activation_io_out_6;
  wire Activation_io_out_5;
  wire Activation_io_out_4;
  wire Activation_io_out_3;
  wire Activation_io_out_2;
  wire Activation_io_out_1;
  wire Activation_io_out_0;
  wire control_io_ready;
  wire control_io_valid;
  wire control_io_done;
  wire[3:0] control_io_selectX;
  wire control_io_memoryRestart;
  wire control_io_chainRestart;
  wire[9:0] Chain_io_ys_9;
  wire[9:0] Chain_io_ys_8;
  wire[9:0] Chain_io_ys_7;
  wire[9:0] Chain_io_ys_6;
  wire[9:0] Chain_io_ys_5;
  wire[9:0] Chain_io_ys_4;
  wire[9:0] Chain_io_ys_3;
  wire[9:0] Chain_io_ys_2;
  wire[9:0] Chain_io_ys_1;
  wire[9:0] Chain_io_ys_0;
  wire[15:0] memoryStreamer_io_weights_9;
  wire[15:0] memoryStreamer_io_weights_8;
  wire[15:0] memoryStreamer_io_weights_7;
  wire[15:0] memoryStreamer_io_weights_6;
  wire[15:0] memoryStreamer_io_weights_5;
  wire[15:0] memoryStreamer_io_weights_4;
  wire[15:0] memoryStreamer_io_weights_3;
  wire[15:0] memoryStreamer_io_weights_2;
  wire[15:0] memoryStreamer_io_weights_1;
  wire[15:0] memoryStreamer_io_weights_0;
  wire[7:0] memoryStreamer_io_bias;


  assign T39 = T0[9:0];
  assign T0 = T1;
  assign T1 = {1'h0, Chain_io_ys_0};
  assign T40 = T2[9:0];
  assign T2 = T3;
  assign T3 = {1'h0, Chain_io_ys_1};
  assign T41 = T4[9:0];
  assign T4 = T5;
  assign T5 = {1'h0, Chain_io_ys_2};
  assign T42 = T6[9:0];
  assign T6 = T7;
  assign T7 = {1'h0, Chain_io_ys_3};
  assign T43 = T8[9:0];
  assign T8 = T9;
  assign T9 = {1'h0, Chain_io_ys_4};
  assign T44 = T10[9:0];
  assign T10 = T11;
  assign T11 = {1'h0, Chain_io_ys_5};
  assign T45 = T12[9:0];
  assign T12 = T13;
  assign T13 = {1'h0, Chain_io_ys_6};
  assign T46 = T14[9:0];
  assign T14 = T15;
  assign T15 = {1'h0, Chain_io_ys_7};
  assign T47 = T16[9:0];
  assign T16 = T17;
  assign T17 = {1'h0, Chain_io_ys_8};
  assign T48 = T18[9:0];
  assign T18 = T19;
  assign T19 = {1'h0, Chain_io_ys_9};
  assign io_done = control_io_done;
  assign io_xOutValid = control_io_valid;
  assign io_xOut_0 = T20;
  assign T20 = T38 ? T36 : T21;
  assign T21 = T35 ? T29 : T22;
  assign T22 = T28 ? T26 : T23;
  assign T23 = T24 ? Activation_io_out_1 : Activation_io_out_0;
  assign T24 = T25[0];
  assign T25 = control_io_selectX;
  assign T26 = T27 ? Activation_io_out_3 : Activation_io_out_2;
  assign T27 = T25[0];
  assign T28 = T25[1];
  assign T29 = T34 ? T32 : T30;
  assign T30 = T31 ? Activation_io_out_5 : Activation_io_out_4;
  assign T31 = T25[0];
  assign T32 = T33 ? Activation_io_out_7 : Activation_io_out_6;
  assign T33 = T25[0];
  assign T34 = T25[1];
  assign T35 = T25[2];
  assign T36 = T37 ? Activation_io_out_9 : Activation_io_out_8;
  assign T37 = T25[0];
  assign T38 = T25[3];
  assign io_startOut = io_start;
  assign io_ready = control_io_ready;
  WarpControl_2 control(.clk(clk), .reset(reset),
       .io_ready( control_io_ready ),
       .io_start( io_start ),
       .io_nextReady( io_pipeReady ),
       .io_valid( control_io_valid ),
       .io_done( control_io_done ),
       .io_selectX( control_io_selectX ),
       .io_memoryRestart( control_io_memoryRestart ),
       .io_chainRestart( control_io_chainRestart )
  );
  Chain_2 Chain(.clk(clk), .reset(reset),
       .io_weights_9( memoryStreamer_io_weights_9 ),
       .io_weights_8( memoryStreamer_io_weights_8 ),
       .io_weights_7( memoryStreamer_io_weights_7 ),
       .io_weights_6( memoryStreamer_io_weights_6 ),
       .io_weights_5( memoryStreamer_io_weights_5 ),
       .io_weights_4( memoryStreamer_io_weights_4 ),
       .io_weights_3( memoryStreamer_io_weights_3 ),
       .io_weights_2( memoryStreamer_io_weights_2 ),
       .io_weights_1( memoryStreamer_io_weights_1 ),
       .io_weights_0( memoryStreamer_io_weights_0 ),
       .io_bias( memoryStreamer_io_bias ),
       .io_restartIn( control_io_chainRestart ),
       .io_xs( io_xIn_0 ),
       .io_ys_9( Chain_io_ys_9 ),
       .io_ys_8( Chain_io_ys_8 ),
       .io_ys_7( Chain_io_ys_7 ),
       .io_ys_6( Chain_io_ys_6 ),
       .io_ys_5( Chain_io_ys_5 ),
       .io_ys_4( Chain_io_ys_4 ),
       .io_ys_3( Chain_io_ys_3 ),
       .io_ys_2( Chain_io_ys_2 ),
       .io_ys_1( Chain_io_ys_1 ),
       .io_ys_0( Chain_io_ys_0 )
  );
  Activation_2 Activation(
       .io_in_9( T48 ),
       .io_in_8( T47 ),
       .io_in_7( T46 ),
       .io_in_6( T45 ),
       .io_in_5( T44 ),
       .io_in_4( T43 ),
       .io_in_3( T42 ),
       .io_in_2( T41 ),
       .io_in_1( T40 ),
       .io_in_0( T39 ),
       .io_out_9( Activation_io_out_9 ),
       .io_out_8( Activation_io_out_8 ),
       .io_out_7( Activation_io_out_7 ),
       .io_out_6( Activation_io_out_6 ),
       .io_out_5( Activation_io_out_5 ),
       .io_out_4( Activation_io_out_4 ),
       .io_out_3( Activation_io_out_3 ),
       .io_out_2( Activation_io_out_2 ),
       .io_out_1( Activation_io_out_1 ),
       .io_out_0( Activation_io_out_0 )
  );
  MemoryStreamer_3 memoryStreamer(.clk(clk), .reset(reset),
       .io_restart( control_io_memoryRestart ),
       .io_weights_9( memoryStreamer_io_weights_9 ),
       .io_weights_8( memoryStreamer_io_weights_8 ),
       .io_weights_7( memoryStreamer_io_weights_7 ),
       .io_weights_6( memoryStreamer_io_weights_6 ),
       .io_weights_5( memoryStreamer_io_weights_5 ),
       .io_weights_4( memoryStreamer_io_weights_4 ),
       .io_weights_3( memoryStreamer_io_weights_3 ),
       .io_weights_2( memoryStreamer_io_weights_2 ),
       .io_weights_1( memoryStreamer_io_weights_1 ),
       .io_weights_0( memoryStreamer_io_weights_0 ),
       .io_bias( memoryStreamer_io_bias )
  );
endmodule

module BitToWord_1(input clk,
    input  io_enable,
    input  io_bit,
    output[15:0] io_word
);

  wire[15:0] T0;
  reg  R1;
  wire T2;
  reg  R3;
  wire T4;
  reg  R5;
  wire T6;
  reg  R7;
  wire T8;
  reg  R9;
  wire T10;
  reg  R11;
  wire T12;
  reg  R13;
  wire T14;
  reg  R15;
  wire T16;
  reg  R17;
  wire T18;
  reg  R19;
  wire T20;
  reg  R21;
  wire T22;
  reg  R23;
  wire T24;
  reg  R25;
  wire T26;
  reg  R27;
  wire T28;
  reg  R29;
  wire T30;
  reg  R31;
  wire T32;
  wire[14:0] T33;
  wire[13:0] T34;
  wire[12:0] T35;
  wire[11:0] T36;
  wire[10:0] T37;
  wire[9:0] T38;
  wire[8:0] T39;
  wire[7:0] T40;
  wire[6:0] T41;
  wire[5:0] T42;
  wire[4:0] T43;
  wire[3:0] T44;
  wire[2:0] T45;
  wire[1:0] T46;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R3 = {1{$random}};
    R5 = {1{$random}};
    R7 = {1{$random}};
    R9 = {1{$random}};
    R11 = {1{$random}};
    R13 = {1{$random}};
    R15 = {1{$random}};
    R17 = {1{$random}};
    R19 = {1{$random}};
    R21 = {1{$random}};
    R23 = {1{$random}};
    R25 = {1{$random}};
    R27 = {1{$random}};
    R29 = {1{$random}};
    R31 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_word = T0;
  assign T0 = {T33, R1};
  assign T2 = io_enable ? R3 : R1;
  assign T4 = io_enable ? R5 : R3;
  assign T6 = io_enable ? R7 : R5;
  assign T8 = io_enable ? R9 : R7;
  assign T10 = io_enable ? R11 : R9;
  assign T12 = io_enable ? R13 : R11;
  assign T14 = io_enable ? R15 : R13;
  assign T16 = io_enable ? R17 : R15;
  assign T18 = io_enable ? R19 : R17;
  assign T20 = io_enable ? R21 : R19;
  assign T22 = io_enable ? R23 : R21;
  assign T24 = io_enable ? R25 : R23;
  assign T26 = io_enable ? R27 : R25;
  assign T28 = io_enable ? R29 : R27;
  assign T30 = io_enable ? R31 : R29;
  assign T32 = io_enable ? io_bit : R31;
  assign T33 = {T34, R3};
  assign T34 = {T35, R5};
  assign T35 = {T36, R7};
  assign T36 = {T37, R9};
  assign T37 = {T38, R11};
  assign T38 = {T39, R13};
  assign T39 = {T40, R15};
  assign T40 = {T41, R17};
  assign T41 = {T42, R19};
  assign T42 = {T43, R21};
  assign T43 = {T44, R23};
  assign T44 = {T45, R25};
  assign T45 = {T46, R27};
  assign T46 = {R31, R29};

  always @(posedge clk) begin
    if(io_enable) begin
      R1 <= R3;
    end
    if(io_enable) begin
      R3 <= R5;
    end
    if(io_enable) begin
      R5 <= R7;
    end
    if(io_enable) begin
      R7 <= R9;
    end
    if(io_enable) begin
      R9 <= R11;
    end
    if(io_enable) begin
      R11 <= R13;
    end
    if(io_enable) begin
      R13 <= R15;
    end
    if(io_enable) begin
      R15 <= R17;
    end
    if(io_enable) begin
      R17 <= R19;
    end
    if(io_enable) begin
      R19 <= R21;
    end
    if(io_enable) begin
      R21 <= R23;
    end
    if(io_enable) begin
      R23 <= R25;
    end
    if(io_enable) begin
      R25 <= R27;
    end
    if(io_enable) begin
      R27 <= R29;
    end
    if(io_enable) begin
      R29 <= R31;
    end
    if(io_enable) begin
      R31 <= io_bit;
    end
  end
endmodule

module AsyncUpDownCounter_0(input clk, input reset,
    input  io_up,
    input  io_down,
    output[3:0] io_value
);

  wire[3:0] T0;
  wire[3:0] T1;
  wire[3:0] T2;
  wire[3:0] T3;
  wire T4;
  wire[3:0] T5;
  wire T6;
  wire T7;
  reg [3:0] reg_;
  wire[3:0] T18;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    reg_ = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = T0;
  assign T0 = T16 ? reg_ : T1;
  assign T1 = T6 ? T5 : T2;
  assign T2 = T4 ? T3 : reg_;
  assign T3 = reg_ + 4'h4;
  assign T4 = io_up & io_down;
  assign T5 = reg_ + 4'h4;
  assign T6 = T7 & io_up;
  assign T7 = T4 ^ 1'h1;
  assign T18 = reset ? 4'h0 : T8;
  assign T8 = T13 ? reg_ : T9;
  assign T9 = T16 ? T12 : T10;
  assign T10 = T6 ? T5 : T11;
  assign T11 = T4 ? reg_ : reg_;
  assign T12 = reg_ - 4'h4;
  assign T13 = T14 ^ 1'h1;
  assign T14 = T15 | io_down;
  assign T15 = T4 | io_up;
  assign T16 = T17 & io_down;
  assign T17 = T15 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      reg_ <= 4'h0;
    end else if(T13) begin
      reg_ <= reg_;
    end else if(T16) begin
      reg_ <= T12;
    end else if(T6) begin
      reg_ <= T5;
    end else if(T4) begin
      reg_ <= reg_;
    end
  end
endmodule

module UpDownCounter_1(input clk, input reset,
    input  io_up,
    input  io_down,
    output[3:0] io_value
);

  reg [3:0] reg_;
  wire[3:0] T10;
  wire[3:0] T0;
  wire[3:0] T1;
  wire[3:0] T2;
  wire T3;
  wire T4;
  wire T5;
  wire[3:0] T6;
  wire T7;
  wire T8;
  wire T9;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    reg_ = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = reg_;
  assign T10 = reset ? 4'h0 : T0;
  assign T0 = T7 ? T6 : T1;
  assign T1 = T3 ? T2 : reg_;
  assign T2 = reg_ + 4'h4;
  assign T3 = T4 & io_up;
  assign T4 = T5 ^ 1'h1;
  assign T5 = io_up & io_down;
  assign T6 = reg_ - 4'h3;
  assign T7 = T8 & io_down;
  assign T8 = T9 ^ 1'h1;
  assign T9 = T5 | io_up;

  always @(posedge clk) begin
    if(reset) begin
      reg_ <= 4'h0;
    end else if(T7) begin
      reg_ <= T6;
    end else if(T3) begin
      reg_ <= T2;
    end
  end
endmodule

module AsyncCounter_1(input clk, input reset,
    input  io_enable,
    output[5:0] io_value
);

  wire[5:0] T0;
  reg [5:0] v;
  wire[5:0] T5;
  wire[5:0] T1;
  wire[5:0] T2;
  wire[5:0] T3;
  wire T4;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    v = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = T0;
  assign T0 = io_enable ? T2 : v;
  assign T5 = reset ? 6'h0 : T1;
  assign T1 = io_enable ? T2 : v;
  assign T2 = T4 ? 6'h0 : T3;
  assign T3 = v + 6'h10;
  assign T4 = v == 6'h20;

  always @(posedge clk) begin
    if(reset) begin
      v <= 6'h0;
    end else if(io_enable) begin
      v <= T2;
    end
  end
endmodule

module CounterWithSyncAndAsyncReset_1(input clk, input reset,
    input  io_enable,
    input  io_syncRst,
    input  io_asyncRst,
    output[3:0] io_value
);

  wire[3:0] T0;
  reg [3:0] v;
  wire[3:0] T13;
  wire[3:0] T1;
  wire[3:0] T2;
  wire[3:0] T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire[3:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire[3:0] T12;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    v = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = T0;
  assign T0 = io_enable ? T12 : v;
  assign T13 = reset ? 4'h0 : T1;
  assign T1 = T9 ? T8 : T2;
  assign T2 = T5 ? 4'h0 : T3;
  assign T3 = T4 ? 4'h1 : v;
  assign T4 = io_enable & io_asyncRst;
  assign T5 = io_enable & T6;
  assign T6 = T7 & io_syncRst;
  assign T7 = io_asyncRst ^ 1'h1;
  assign T8 = v + 4'h1;
  assign T9 = io_enable & T10;
  assign T10 = T11 ^ 1'h1;
  assign T11 = io_asyncRst | io_syncRst;
  assign T12 = io_asyncRst ? 4'h0 : v;

  always @(posedge clk) begin
    if(reset) begin
      v <= 4'h0;
    end else if(T9) begin
      v <= T8;
    end else if(T5) begin
      v <= 4'h0;
    end else if(T4) begin
      v <= 4'h1;
    end
  end
endmodule

module CircularPeekQueue_1(input clk, input reset,
    input  io_writeEnable,
    input  io_nextBlock,
    input [15:0] io_input,
    output[15:0] io_output
);

  reg [5:0] writeAddr;
  wire[5:0] T10;
  wire[5:0] T0;
  wire[5:0] T1;
  wire T2;
  wire T3;
  wire[5:0] T4;
  wire T5;
  wire T6;
  wire[5:0] T7;
  wire[5:0] T11;
  wire[3:0] T8;
  wire T9;
  wire[5:0] currentBlockOffset_io_value;
  wire[3:0] inBlockReadOffset_io_value;
  wire[15:0] queue_b_dout;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    writeAddr = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T10 = reset ? 6'h10 : T0;
  assign T0 = T5 ? T4 : T1;
  assign T1 = T2 ? 6'h0 : writeAddr;
  assign T2 = io_writeEnable & T3;
  assign T3 = writeAddr == 6'h2f;
  assign T4 = writeAddr + 6'h1;
  assign T5 = io_writeEnable & T6;
  assign T6 = T3 ^ 1'h1;
  assign T7 = currentBlockOffset_io_value + T11;
  assign T11 = {2'h0, T8};
  assign T8 = io_nextBlock ? 4'h0 : inBlockReadOffset_io_value;
  assign T9 = inBlockReadOffset_io_value == 4'hf;
  assign io_output = queue_b_dout;
  AsyncCounter_1 currentBlockOffset(.clk(clk), .reset(reset),
       .io_enable( io_nextBlock ),
       .io_value( currentBlockOffset_io_value )
  );
  CounterWithSyncAndAsyncReset_1 inBlockReadOffset(.clk(clk), .reset(reset),
       .io_enable( 1'h1 ),
       .io_syncRst( T9 ),
       .io_asyncRst( io_nextBlock ),
       .io_value( inBlockReadOffset_io_value )
  );
  DualPortBRAM # (
    .DATA(16),
    .ADDR(6)
  ) queue(.clk(clk),
       .b_addr( T7 ),
       //.b_din(  )
       .b_wr( 1'h0 ),
       .b_dout( queue_b_dout ),
       .a_addr( writeAddr ),
       .a_din( io_input ),
       .a_wr( io_writeEnable )
       //.a_dout(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign queue.b_din = {1{$random}};
// synthesis translate_on
`endif

  always @(posedge clk) begin
    if(reset) begin
      writeAddr <= 6'h10;
    end else if(T5) begin
      writeAddr <= T4;
    end else if(T2) begin
      writeAddr <= 6'h0;
    end
  end
endmodule

module WrappingCounter_0(
    input  io_enable,
    output io_value
);



  assign io_value = 1'h0;
endmodule

module WrappingCounter_1(
    input  io_enable,
    output io_value
);



  assign io_value = 1'h1;
endmodule

module WrappingCounter_2(
    input  io_enable,
    output[1:0] io_value
);



  assign io_value = 2'h2;
endmodule

module WrappingCounter_3(
    input  io_enable,
    output[1:0] io_value
);



  assign io_value = 2'h3;
endmodule

module WrappingCounter_4(input clk, input reset,
    input  io_enable,
    output[2:0] io_value
);

  reg [2:0] R0;
  wire[2:0] T11;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire T5;
  wire T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire T9;
  wire T10;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = R0;
  assign T11 = reset ? 3'h1 : T1;
  assign T1 = T9 ? T8 : T2;
  assign T2 = T5 ? T3 : R0;
  assign T3 = T4 - 3'h4;
  assign T4 = R0 + 3'h3;
  assign T5 = io_enable & T6;
  assign T6 = 3'h4 <= T7;
  assign T7 = R0 + 3'h3;
  assign T8 = R0 + 3'h3;
  assign T9 = io_enable & T10;
  assign T10 = T6 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R0 <= 3'h1;
    end else if(T9) begin
      R0 <= T8;
    end else if(T5) begin
      R0 <= T3;
    end
  end
endmodule

module WrappingCounter_5(input clk, input reset,
    input  io_enable,
    output[2:0] io_value
);

  reg [2:0] R0;
  wire[2:0] T11;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire T5;
  wire T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire T9;
  wire T10;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = R0;
  assign T11 = reset ? 3'h2 : T1;
  assign T1 = T9 ? T8 : T2;
  assign T2 = T5 ? T3 : R0;
  assign T3 = T4 - 3'h4;
  assign T4 = R0 + 3'h3;
  assign T5 = io_enable & T6;
  assign T6 = 3'h4 <= T7;
  assign T7 = R0 + 3'h3;
  assign T8 = R0 + 3'h3;
  assign T9 = io_enable & T10;
  assign T10 = T6 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R0 <= 3'h2;
    end else if(T9) begin
      R0 <= T8;
    end else if(T5) begin
      R0 <= T3;
    end
  end
endmodule

module WrappingCounter_6(input clk, input reset,
    input  io_enable,
    output[2:0] io_value
);

  reg [2:0] R0;
  wire[2:0] T11;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire T5;
  wire T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire T9;
  wire T10;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = R0;
  assign T11 = reset ? 3'h3 : T1;
  assign T1 = T9 ? T8 : T2;
  assign T2 = T5 ? T3 : R0;
  assign T3 = T4 - 3'h4;
  assign T4 = R0 + 3'h3;
  assign T5 = io_enable & T6;
  assign T6 = 3'h4 <= T7;
  assign T7 = R0 + 3'h3;
  assign T8 = R0 + 3'h3;
  assign T9 = io_enable & T10;
  assign T10 = T6 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R0 <= 3'h3;
    end else if(T9) begin
      R0 <= T8;
    end else if(T5) begin
      R0 <= T3;
    end
  end
endmodule

module WrappingCounter_7(input clk, input reset,
    input  io_enable,
    output[2:0] io_value
);

  reg [2:0] R0;
  wire[2:0] T11;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire T5;
  wire T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire T9;
  wire T10;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = R0;
  assign T11 = reset ? 3'h0 : T1;
  assign T1 = T9 ? T8 : T2;
  assign T2 = T5 ? T3 : R0;
  assign T3 = T4 - 3'h4;
  assign T4 = R0 + 3'h1;
  assign T5 = io_enable & T6;
  assign T6 = 3'h4 <= T7;
  assign T7 = R0 + 3'h1;
  assign T8 = R0 + 3'h1;
  assign T9 = io_enable & T10;
  assign T10 = T6 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R0 <= 3'h0;
    end else if(T9) begin
      R0 <= T8;
    end else if(T5) begin
      R0 <= T3;
    end
  end
endmodule

module WrappingCounter_8(input clk, input reset,
    input  io_enable,
    output[2:0] io_value
);

  reg [2:0] R0;
  wire[2:0] T11;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire T5;
  wire T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire T9;
  wire T10;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = R0;
  assign T11 = reset ? 3'h1 : T1;
  assign T1 = T9 ? T8 : T2;
  assign T2 = T5 ? T3 : R0;
  assign T3 = T4 - 3'h4;
  assign T4 = R0 + 3'h1;
  assign T5 = io_enable & T6;
  assign T6 = 3'h4 <= T7;
  assign T7 = R0 + 3'h1;
  assign T8 = R0 + 3'h1;
  assign T9 = io_enable & T10;
  assign T10 = T6 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R0 <= 3'h1;
    end else if(T9) begin
      R0 <= T8;
    end else if(T5) begin
      R0 <= T3;
    end
  end
endmodule

module WrappingCounter_9(input clk, input reset,
    input  io_enable,
    output[2:0] io_value
);

  reg [2:0] R0;
  wire[2:0] T11;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire T5;
  wire T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire T9;
  wire T10;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = R0;
  assign T11 = reset ? 3'h2 : T1;
  assign T1 = T9 ? T8 : T2;
  assign T2 = T5 ? T3 : R0;
  assign T3 = T4 - 3'h4;
  assign T4 = R0 + 3'h1;
  assign T5 = io_enable & T6;
  assign T6 = 3'h4 <= T7;
  assign T7 = R0 + 3'h1;
  assign T8 = R0 + 3'h1;
  assign T9 = io_enable & T10;
  assign T10 = T6 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R0 <= 3'h2;
    end else if(T9) begin
      R0 <= T8;
    end else if(T5) begin
      R0 <= T3;
    end
  end
endmodule

module WrappingCounter_10(input clk, input reset,
    input  io_enable,
    output[2:0] io_value
);

  reg [2:0] R0;
  wire[2:0] T11;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire T5;
  wire T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire T9;
  wire T10;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = R0;
  assign T11 = reset ? 3'h3 : T1;
  assign T1 = T9 ? T8 : T2;
  assign T2 = T5 ? T3 : R0;
  assign T3 = T4 - 3'h4;
  assign T4 = R0 + 3'h1;
  assign T5 = io_enable & T6;
  assign T6 = 3'h4 <= T7;
  assign T7 = R0 + 3'h1;
  assign T8 = R0 + 3'h1;
  assign T9 = io_enable & T10;
  assign T10 = T6 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R0 <= 3'h3;
    end else if(T9) begin
      R0 <= T8;
    end else if(T5) begin
      R0 <= T3;
    end
  end
endmodule

module GearBox_0(input clk, input reset,
    input  io_xsIn_3,
    input  io_xsIn_2,
    input  io_xsIn_1,
    input  io_xsIn_0,
    input  io_validIn,
    input  io_prevDone,
    input  io_prevStart,
    output io_ready,
    input  io_nextReady,
    output io_startNext,
    output[15:0] io_xsOut_2,
    output[15:0] io_xsOut_1,
    output[15:0] io_xsOut_0
);

  wire signalNewPeekBlock;
  wire T0;
  reg  R1;
  wire T76;
  reg  R2;
  wire T77;
  reg  R3;
  wire T78;
  reg  R4;
  wire T79;
  wire[15:0] T5;
  wire[15:0] T6;
  wire T7;
  wire[1:0] T8;
  wire[15:0] T9;
  wire T10;
  wire T11;
  wire T12;
  reg  T13;
  wire[1:0] T80;
  wire T15;
  reg  T16;
  reg  signalBitBuffersFull;
  wire T81;
  wire T18;
  wire signalResetBitBuffers;
  wire[15:0] T19;
  wire[15:0] T20;
  wire T21;
  wire[1:0] T22;
  wire[15:0] T23;
  wire T24;
  wire T25;
  wire T26;
  reg  T27;
  wire[1:0] T82;
  wire T28;
  reg  T29;
  wire[15:0] T30;
  wire[15:0] T31;
  wire T32;
  wire[1:0] T33;
  wire[1:0] T83;
  wire[15:0] T34;
  wire T35;
  wire T36;
  wire T37;
  reg  T38;
  wire[1:0] T84;
  wire T39;
  reg  T40;
  wire[1:0] T85;
  wire[15:0] T41;
  wire[15:0] T42;
  wire T43;
  wire[1:0] T44;
  wire[1:0] T86;
  wire[15:0] T45;
  wire T46;
  wire T47;
  wire T48;
  reg  T49;
  wire[1:0] T87;
  wire T50;
  reg  T51;
  wire[1:0] T88;
  reg  R52;
  wire T89;
  reg  R53;
  wire T90;
  wire[15:0] T54;
  wire[15:0] T55;
  wire T56;
  wire[1:0] T57;
  wire[1:0] T91;
  wire[15:0] T58;
  wire T59;
  wire T60;
  wire[15:0] T61;
  wire[15:0] T62;
  wire T63;
  wire[1:0] T64;
  wire[1:0] T92;
  wire[15:0] T65;
  wire T66;
  wire T67;
  wire[15:0] T68;
  wire[15:0] T69;
  wire T70;
  wire[1:0] T71;
  wire[1:0] T93;
  wire[15:0] T72;
  wire T73;
  wire T74;
  reg  R75;
  wire T94;
  wire hasEnoughEmptyBlocks;
  wire[3:0] reservedBlocks;
  wire[15:0] BitToWord_io_word;
  wire[15:0] BitToWord_1_io_word;
  wire[15:0] BitToWord_2_io_word;
  wire[15:0] BitToWord_3_io_word;
  wire[3:0] fillingBlock_io_value;
  wire[3:0] bitCounter_io_value;
  wire[3:0] blocksReady_io_value;
  wire inputSelectCounter_io_value;
  wire inputSelectCounter_1_io_value;
  wire[1:0] inputSelectCounter_2_io_value;
  wire[1:0] inputSelectCounter_3_io_value;
  wire[2:0] queueOutputSelectCounters_io_value;
  wire[2:0] queueOutputSelectCounters_1_io_value;
  wire[2:0] queueOutputSelectCounters_2_io_value;
  wire[2:0] outputSelectCounters_io_value;
  wire[2:0] outputSelectCounters_1_io_value;
  wire[2:0] outputSelectCounters_2_io_value;
  wire[2:0] outputSelectCounters_3_io_value;
  wire[15:0] CircularPeekQueue_io_output;
  wire[15:0] CircularPeekQueue_1_io_output;
  wire[15:0] CircularPeekQueue_2_io_output;
  wire[15:0] CircularPeekQueue_3_io_output;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R2 = {1{$random}};
    R3 = {1{$random}};
    R4 = {1{$random}};
    signalBitBuffersFull = {1{$random}};
    R52 = {1{$random}};
    R53 = {1{$random}};
    R75 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign signalNewPeekBlock = io_nextReady & T0;
  assign T0 = 4'h3 <= blocksReady_io_value;
  assign T76 = reset ? 1'h0 : io_prevDone;
  assign T77 = reset ? 1'h0 : io_prevDone;
  assign T78 = reset ? 1'h0 : io_prevDone;
  assign T79 = reset ? 1'h0 : io_prevDone;
  assign T5 = T11 ? T9 : T6;
  assign T6 = T7 ? BitToWord_1_io_word : BitToWord_io_word;
  assign T7 = T8[0];
  assign T8 = inputSelectCounter_3_io_value;
  assign T9 = T10 ? BitToWord_3_io_word : BitToWord_2_io_word;
  assign T10 = T8[0];
  assign T11 = T8[1];
  assign T12 = signalNewPeekBlock & T13;
  always @(*) case (T80)
    0: T13 = 1'h1;
    1: T13 = 1'h1;
    2: T13 = 1'h1;
    3: T13 = 1'h0;
    default: begin
      T13 = 1'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T13 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T80 = outputSelectCounters_3_io_value[1:0];
  assign T15 = signalBitBuffersFull & T16;
  always @(*) case (inputSelectCounter_3_io_value)
    0: T16 = 1'h1;
    1: T16 = 1'h1;
    2: T16 = 1'h1;
    3: T16 = 1'h1;
    default: begin
      T16 = 1'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T16 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T81 = reset ? 1'h0 : T18;
  assign T18 = io_validIn & signalResetBitBuffers;
  assign signalResetBitBuffers = bitCounter_io_value == 4'hf;
  assign T19 = T25 ? T23 : T20;
  assign T20 = T21 ? BitToWord_1_io_word : BitToWord_io_word;
  assign T21 = T22[0];
  assign T22 = inputSelectCounter_2_io_value;
  assign T23 = T24 ? BitToWord_3_io_word : BitToWord_2_io_word;
  assign T24 = T22[0];
  assign T25 = T22[1];
  assign T26 = signalNewPeekBlock & T27;
  always @(*) case (T82)
    0: T27 = 1'h1;
    1: T27 = 1'h1;
    2: T27 = 1'h1;
    3: T27 = 1'h0;
    default: begin
      T27 = 1'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T27 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T82 = outputSelectCounters_2_io_value[1:0];
  assign T28 = signalBitBuffersFull & T29;
  always @(*) case (inputSelectCounter_2_io_value)
    0: T29 = 1'h1;
    1: T29 = 1'h1;
    2: T29 = 1'h1;
    3: T29 = 1'h1;
    default: begin
      T29 = 1'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T29 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T30 = T36 ? T34 : T31;
  assign T31 = T32 ? BitToWord_1_io_word : BitToWord_io_word;
  assign T32 = T33[0];
  assign T33 = T83;
  assign T83 = {1'h0, inputSelectCounter_1_io_value};
  assign T34 = T35 ? BitToWord_3_io_word : BitToWord_2_io_word;
  assign T35 = T33[0];
  assign T36 = T33[1];
  assign T37 = signalNewPeekBlock & T38;
  always @(*) case (T84)
    0: T38 = 1'h1;
    1: T38 = 1'h1;
    2: T38 = 1'h1;
    3: T38 = 1'h0;
    default: begin
      T38 = 1'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T38 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T84 = outputSelectCounters_1_io_value[1:0];
  assign T39 = signalBitBuffersFull & T40;
  always @(*) case (T85)
    0: T40 = 1'h1;
    1: T40 = 1'h1;
    2: T40 = 1'h1;
    3: T40 = 1'h1;
    default: begin
      T40 = 1'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T40 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T85 = {1'h0, inputSelectCounter_1_io_value};
  assign T41 = T47 ? T45 : T42;
  assign T42 = T43 ? BitToWord_1_io_word : BitToWord_io_word;
  assign T43 = T44[0];
  assign T44 = T86;
  assign T86 = {1'h0, inputSelectCounter_io_value};
  assign T45 = T46 ? BitToWord_3_io_word : BitToWord_2_io_word;
  assign T46 = T44[0];
  assign T47 = T44[1];
  assign T48 = signalNewPeekBlock & T49;
  always @(*) case (T87)
    0: T49 = 1'h1;
    1: T49 = 1'h1;
    2: T49 = 1'h1;
    3: T49 = 1'h0;
    default: begin
      T49 = 1'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T49 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T87 = outputSelectCounters_io_value[1:0];
  assign T50 = signalBitBuffersFull & T51;
  always @(*) case (T88)
    0: T51 = 1'h1;
    1: T51 = 1'h1;
    2: T51 = 1'h1;
    3: T51 = 1'h1;
    default: begin
      T51 = 1'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T51 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T88 = {1'h0, inputSelectCounter_io_value};
  assign T89 = reset ? 1'h0 : io_prevDone;
  assign T90 = reset ? 1'h0 : io_prevDone;
  assign io_xsOut_0 = T54;
  assign T54 = T60 ? T58 : T55;
  assign T55 = T56 ? CircularPeekQueue_1_io_output : CircularPeekQueue_io_output;
  assign T56 = T57[0];
  assign T57 = T91;
  assign T91 = queueOutputSelectCounters_io_value[1:0];
  assign T58 = T59 ? CircularPeekQueue_3_io_output : CircularPeekQueue_2_io_output;
  assign T59 = T57[0];
  assign T60 = T57[1];
  assign io_xsOut_1 = T61;
  assign T61 = T67 ? T65 : T62;
  assign T62 = T63 ? CircularPeekQueue_1_io_output : CircularPeekQueue_io_output;
  assign T63 = T64[0];
  assign T64 = T92;
  assign T92 = queueOutputSelectCounters_1_io_value[1:0];
  assign T65 = T66 ? CircularPeekQueue_3_io_output : CircularPeekQueue_2_io_output;
  assign T66 = T64[0];
  assign T67 = T64[1];
  assign io_xsOut_2 = T68;
  assign T68 = T74 ? T72 : T69;
  assign T69 = T70 ? CircularPeekQueue_1_io_output : CircularPeekQueue_io_output;
  assign T70 = T71[0];
  assign T71 = T93;
  assign T93 = queueOutputSelectCounters_2_io_value[1:0];
  assign T72 = T73 ? CircularPeekQueue_3_io_output : CircularPeekQueue_2_io_output;
  assign T73 = T71[0];
  assign T74 = T71[1];
  assign io_startNext = R75;
  assign T94 = reset ? 1'h0 : signalNewPeekBlock;
  assign io_ready = hasEnoughEmptyBlocks;
  assign hasEnoughEmptyBlocks = reservedBlocks <= 4'h5;
  assign reservedBlocks = blocksReady_io_value + fillingBlock_io_value;
  BitToWord_1 BitToWord(.clk(clk),
       .io_enable( io_validIn ),
       .io_bit( io_xsIn_0 ),
       .io_word( BitToWord_io_word )
  );
  BitToWord_1 BitToWord_1(.clk(clk),
       .io_enable( io_validIn ),
       .io_bit( io_xsIn_1 ),
       .io_word( BitToWord_1_io_word )
  );
  BitToWord_1 BitToWord_2(.clk(clk),
       .io_enable( io_validIn ),
       .io_bit( io_xsIn_2 ),
       .io_word( BitToWord_2_io_word )
  );
  BitToWord_1 BitToWord_3(.clk(clk),
       .io_enable( io_validIn ),
       .io_bit( io_xsIn_3 ),
       .io_word( BitToWord_3_io_word )
  );
  AsyncUpDownCounter_0 fillingBlock(.clk(clk), .reset(reset),
       .io_up( io_prevStart ),
       .io_down( R53 ),
       .io_value( fillingBlock_io_value )
  );
  Counter_2 bitCounter(.clk(clk), .reset(reset),
       .io_enable( io_validIn ),
       .io_rst( signalResetBitBuffers ),
       .io_value( bitCounter_io_value )
  );
  UpDownCounter_1 blocksReady(.clk(clk), .reset(reset),
       .io_up( R52 ),
       .io_down( signalNewPeekBlock ),
       .io_value( blocksReady_io_value )
  );
  CircularPeekQueue_1 CircularPeekQueue(.clk(clk), .reset(reset),
       .io_writeEnable( T50 ),
       .io_nextBlock( T48 ),
       .io_input( T41 ),
       .io_output( CircularPeekQueue_io_output )
  );
  CircularPeekQueue_1 CircularPeekQueue_1(.clk(clk), .reset(reset),
       .io_writeEnable( T39 ),
       .io_nextBlock( T37 ),
       .io_input( T30 ),
       .io_output( CircularPeekQueue_1_io_output )
  );
  CircularPeekQueue_1 CircularPeekQueue_2(.clk(clk), .reset(reset),
       .io_writeEnable( T28 ),
       .io_nextBlock( T26 ),
       .io_input( T19 ),
       .io_output( CircularPeekQueue_2_io_output )
  );
  CircularPeekQueue_1 CircularPeekQueue_3(.clk(clk), .reset(reset),
       .io_writeEnable( T15 ),
       .io_nextBlock( T12 ),
       .io_input( T5 ),
       .io_output( CircularPeekQueue_3_io_output )
  );
  WrappingCounter_0 inputSelectCounter(
       .io_enable( R4 ),
       .io_value( inputSelectCounter_io_value )
  );
  WrappingCounter_1 inputSelectCounter_1(
       .io_enable( R3 ),
       .io_value( inputSelectCounter_1_io_value )
  );
  WrappingCounter_2 inputSelectCounter_2(
       .io_enable( R2 ),
       .io_value( inputSelectCounter_2_io_value )
  );
  WrappingCounter_3 inputSelectCounter_3(
       .io_enable( R1 ),
       .io_value( inputSelectCounter_3_io_value )
  );
  WrappingCounter_4 queueOutputSelectCounters(.clk(clk), .reset(reset),
       .io_enable( signalNewPeekBlock ),
       .io_value( queueOutputSelectCounters_io_value )
  );
  WrappingCounter_5 queueOutputSelectCounters_1(.clk(clk), .reset(reset),
       .io_enable( signalNewPeekBlock ),
       .io_value( queueOutputSelectCounters_1_io_value )
  );
  WrappingCounter_6 queueOutputSelectCounters_2(.clk(clk), .reset(reset),
       .io_enable( signalNewPeekBlock ),
       .io_value( queueOutputSelectCounters_2_io_value )
  );
  WrappingCounter_7 outputSelectCounters(.clk(clk), .reset(reset),
       .io_enable( signalNewPeekBlock ),
       .io_value( outputSelectCounters_io_value )
  );
  WrappingCounter_8 outputSelectCounters_1(.clk(clk), .reset(reset),
       .io_enable( signalNewPeekBlock ),
       .io_value( outputSelectCounters_1_io_value )
  );
  WrappingCounter_9 outputSelectCounters_2(.clk(clk), .reset(reset),
       .io_enable( signalNewPeekBlock ),
       .io_value( outputSelectCounters_2_io_value )
  );
  WrappingCounter_10 outputSelectCounters_3(.clk(clk), .reset(reset),
       .io_enable( signalNewPeekBlock ),
       .io_value( outputSelectCounters_3_io_value )
  );

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else begin
      R1 <= io_prevDone;
    end
    if(reset) begin
      R2 <= 1'h0;
    end else begin
      R2 <= io_prevDone;
    end
    if(reset) begin
      R3 <= 1'h0;
    end else begin
      R3 <= io_prevDone;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else begin
      R4 <= io_prevDone;
    end
    if(reset) begin
      signalBitBuffersFull <= 1'h0;
    end else begin
      signalBitBuffersFull <= T18;
    end
    if(reset) begin
      R52 <= 1'h0;
    end else begin
      R52 <= io_prevDone;
    end
    if(reset) begin
      R53 <= 1'h0;
    end else begin
      R53 <= io_prevDone;
    end
    if(reset) begin
      R75 <= 1'h0;
    end else begin
      R75 <= signalNewPeekBlock;
    end
  end
endmodule

module AsyncUpDownCounter_1(input clk, input reset,
    input  io_up,
    input  io_down,
    output[2:0] io_value
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire T4;
  wire[2:0] T5;
  wire T6;
  wire T7;
  reg [2:0] reg_;
  wire[2:0] T18;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    reg_ = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = T0;
  assign T0 = T16 ? reg_ : T1;
  assign T1 = T6 ? T5 : T2;
  assign T2 = T4 ? T3 : reg_;
  assign T3 = reg_ + 3'h3;
  assign T4 = io_up & io_down;
  assign T5 = reg_ + 3'h3;
  assign T6 = T7 & io_up;
  assign T7 = T4 ^ 1'h1;
  assign T18 = reset ? 3'h0 : T8;
  assign T8 = T13 ? reg_ : T9;
  assign T9 = T16 ? T12 : T10;
  assign T10 = T6 ? T5 : T11;
  assign T11 = T4 ? reg_ : reg_;
  assign T12 = reg_ - 3'h3;
  assign T13 = T14 ^ 1'h1;
  assign T14 = T15 | io_down;
  assign T15 = T4 | io_up;
  assign T16 = T17 & io_down;
  assign T17 = T15 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      reg_ <= 3'h0;
    end else if(T13) begin
      reg_ <= reg_;
    end else if(T16) begin
      reg_ <= T12;
    end else if(T6) begin
      reg_ <= T5;
    end else if(T4) begin
      reg_ <= reg_;
    end
  end
endmodule

module UpDownCounter_2(input clk, input reset,
    input  io_up,
    input  io_down,
    output[2:0] io_value
);

  reg [2:0] reg_;
  wire[2:0] T10;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire T3;
  wire T4;
  wire T5;
  wire[2:0] T6;
  wire T7;
  wire T8;
  wire T9;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    reg_ = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = reg_;
  assign T10 = reset ? 3'h0 : T0;
  assign T0 = T7 ? T6 : T1;
  assign T1 = T3 ? T2 : reg_;
  assign T2 = reg_ + 3'h3;
  assign T3 = T4 & io_up;
  assign T4 = T5 ^ 1'h1;
  assign T5 = io_up & io_down;
  assign T6 = reg_ - 3'h3;
  assign T7 = T8 & io_down;
  assign T8 = T9 ^ 1'h1;
  assign T9 = T5 | io_up;

  always @(posedge clk) begin
    if(reset) begin
      reg_ <= 3'h0;
    end else if(T7) begin
      reg_ <= T6;
    end else if(T3) begin
      reg_ <= T2;
    end
  end
endmodule

module GearBox_1(input clk, input reset,
    input  io_xsIn_2,
    input  io_xsIn_1,
    input  io_xsIn_0,
    input  io_validIn,
    input  io_prevDone,
    input  io_prevStart,
    output io_ready,
    input  io_nextReady,
    output io_startNext,
    output[15:0] io_xsOut_2,
    output[15:0] io_xsOut_1,
    output[15:0] io_xsOut_0
);

  wire signalNewPeekBlock;
  wire T0;
  reg  R1;
  wire T52;
  reg  R2;
  wire T53;
  reg  R3;
  wire T54;
  wire[15:0] T4;
  wire[15:0] T5;
  wire T6;
  wire[1:0] T7;
  wire T8;
  wire T9;
  reg  T10;
  wire T12;
  reg  T13;
  reg  signalBitBuffersFull;
  wire T55;
  wire T15;
  wire signalResetBitBuffers;
  wire[15:0] T16;
  wire[15:0] T17;
  wire T18;
  wire[1:0] T19;
  wire[1:0] T56;
  wire T20;
  wire T21;
  reg  T22;
  wire[1:0] T57;
  wire T23;
  reg  T24;
  wire[1:0] T58;
  wire[15:0] T25;
  wire[15:0] T26;
  wire T27;
  wire[1:0] T28;
  wire[1:0] T59;
  wire T29;
  wire T30;
  reg  T31;
  wire[1:0] T60;
  wire T32;
  reg  T33;
  wire[1:0] T61;
  reg  R34;
  wire T62;
  reg  R35;
  wire T63;
  wire[15:0] T36;
  wire[15:0] T37;
  wire T38;
  wire[1:0] T39;
  wire[1:0] T64;
  wire T40;
  wire[15:0] T41;
  wire[15:0] T42;
  wire T43;
  wire[1:0] T44;
  wire[1:0] T65;
  wire T45;
  wire[15:0] T46;
  wire[15:0] T47;
  wire T48;
  wire[1:0] T49;
  wire T50;
  reg  R51;
  wire T66;
  wire hasEnoughEmptyBlocks;
  wire[2:0] reservedBlocks;
  wire[15:0] BitToWord_io_word;
  wire[15:0] BitToWord_1_io_word;
  wire[15:0] BitToWord_2_io_word;
  wire[2:0] fillingBlock_io_value;
  wire[3:0] bitCounter_io_value;
  wire[2:0] blocksReady_io_value;
  wire inputSelectCounter_io_value;
  wire inputSelectCounter_1_io_value;
  wire[1:0] inputSelectCounter_2_io_value;
  wire queueOutputSelectCounters_io_value;
  wire queueOutputSelectCounters_1_io_value;
  wire[1:0] queueOutputSelectCounters_2_io_value;
  wire outputSelectCounters_io_value;
  wire outputSelectCounters_1_io_value;
  wire[1:0] outputSelectCounters_2_io_value;
  wire[15:0] CircularPeekQueue_io_output;
  wire[15:0] CircularPeekQueue_1_io_output;
  wire[15:0] CircularPeekQueue_2_io_output;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R2 = {1{$random}};
    R3 = {1{$random}};
    signalBitBuffersFull = {1{$random}};
    R34 = {1{$random}};
    R35 = {1{$random}};
    R51 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign signalNewPeekBlock = io_nextReady & T0;
  assign T0 = 3'h3 <= blocksReady_io_value;
  assign T52 = reset ? 1'h0 : io_prevDone;
  assign T53 = reset ? 1'h0 : io_prevDone;
  assign T54 = reset ? 1'h0 : io_prevDone;
  assign T4 = T8 ? BitToWord_2_io_word : T5;
  assign T5 = T6 ? BitToWord_1_io_word : BitToWord_io_word;
  assign T6 = T7[0];
  assign T7 = inputSelectCounter_2_io_value;
  assign T8 = T7[1];
  assign T9 = signalNewPeekBlock & T10;
  always @(*) case (outputSelectCounters_2_io_value)
    0: T10 = 1'h1;
    1: T10 = 1'h1;
    2: T10 = 1'h1;
    default: begin
      T10 = 1'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T10 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T12 = signalBitBuffersFull & T13;
  always @(*) case (inputSelectCounter_2_io_value)
    0: T13 = 1'h1;
    1: T13 = 1'h1;
    2: T13 = 1'h1;
    default: begin
      T13 = 1'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T13 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T55 = reset ? 1'h0 : T15;
  assign T15 = io_validIn & signalResetBitBuffers;
  assign signalResetBitBuffers = bitCounter_io_value == 4'hf;
  assign T16 = T20 ? BitToWord_2_io_word : T17;
  assign T17 = T18 ? BitToWord_1_io_word : BitToWord_io_word;
  assign T18 = T19[0];
  assign T19 = T56;
  assign T56 = {1'h0, inputSelectCounter_1_io_value};
  assign T20 = T19[1];
  assign T21 = signalNewPeekBlock & T22;
  always @(*) case (T57)
    0: T22 = 1'h1;
    1: T22 = 1'h1;
    2: T22 = 1'h1;
    default: begin
      T22 = 1'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T22 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T57 = {1'h0, outputSelectCounters_1_io_value};
  assign T23 = signalBitBuffersFull & T24;
  always @(*) case (T58)
    0: T24 = 1'h1;
    1: T24 = 1'h1;
    2: T24 = 1'h1;
    default: begin
      T24 = 1'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T24 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T58 = {1'h0, inputSelectCounter_1_io_value};
  assign T25 = T29 ? BitToWord_2_io_word : T26;
  assign T26 = T27 ? BitToWord_1_io_word : BitToWord_io_word;
  assign T27 = T28[0];
  assign T28 = T59;
  assign T59 = {1'h0, inputSelectCounter_io_value};
  assign T29 = T28[1];
  assign T30 = signalNewPeekBlock & T31;
  always @(*) case (T60)
    0: T31 = 1'h1;
    1: T31 = 1'h1;
    2: T31 = 1'h1;
    default: begin
      T31 = 1'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T31 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T60 = {1'h0, outputSelectCounters_io_value};
  assign T32 = signalBitBuffersFull & T33;
  always @(*) case (T61)
    0: T33 = 1'h1;
    1: T33 = 1'h1;
    2: T33 = 1'h1;
    default: begin
      T33 = 1'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T33 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T61 = {1'h0, inputSelectCounter_io_value};
  assign T62 = reset ? 1'h0 : io_prevDone;
  assign T63 = reset ? 1'h0 : io_prevDone;
  assign io_xsOut_0 = T36;
  assign T36 = T40 ? CircularPeekQueue_2_io_output : T37;
  assign T37 = T38 ? CircularPeekQueue_1_io_output : CircularPeekQueue_io_output;
  assign T38 = T39[0];
  assign T39 = T64;
  assign T64 = {1'h0, queueOutputSelectCounters_io_value};
  assign T40 = T39[1];
  assign io_xsOut_1 = T41;
  assign T41 = T45 ? CircularPeekQueue_2_io_output : T42;
  assign T42 = T43 ? CircularPeekQueue_1_io_output : CircularPeekQueue_io_output;
  assign T43 = T44[0];
  assign T44 = T65;
  assign T65 = {1'h0, queueOutputSelectCounters_1_io_value};
  assign T45 = T44[1];
  assign io_xsOut_2 = T46;
  assign T46 = T50 ? CircularPeekQueue_2_io_output : T47;
  assign T47 = T48 ? CircularPeekQueue_1_io_output : CircularPeekQueue_io_output;
  assign T48 = T49[0];
  assign T49 = queueOutputSelectCounters_2_io_value;
  assign T50 = T49[1];
  assign io_startNext = R51;
  assign T66 = reset ? 1'h0 : signalNewPeekBlock;
  assign io_ready = hasEnoughEmptyBlocks;
  assign hasEnoughEmptyBlocks = reservedBlocks <= 3'h3;
  assign reservedBlocks = blocksReady_io_value + fillingBlock_io_value;
  BitToWord_1 BitToWord(.clk(clk),
       .io_enable( io_validIn ),
       .io_bit( io_xsIn_0 ),
       .io_word( BitToWord_io_word )
  );
  BitToWord_1 BitToWord_1(.clk(clk),
       .io_enable( io_validIn ),
       .io_bit( io_xsIn_1 ),
       .io_word( BitToWord_1_io_word )
  );
  BitToWord_1 BitToWord_2(.clk(clk),
       .io_enable( io_validIn ),
       .io_bit( io_xsIn_2 ),
       .io_word( BitToWord_2_io_word )
  );
  AsyncUpDownCounter_1 fillingBlock(.clk(clk), .reset(reset),
       .io_up( io_prevStart ),
       .io_down( R35 ),
       .io_value( fillingBlock_io_value )
  );
  Counter_2 bitCounter(.clk(clk), .reset(reset),
       .io_enable( io_validIn ),
       .io_rst( signalResetBitBuffers ),
       .io_value( bitCounter_io_value )
  );
  UpDownCounter_2 blocksReady(.clk(clk), .reset(reset),
       .io_up( R34 ),
       .io_down( signalNewPeekBlock ),
       .io_value( blocksReady_io_value )
  );
  CircularPeekQueue_1 CircularPeekQueue(.clk(clk), .reset(reset),
       .io_writeEnable( T32 ),
       .io_nextBlock( T30 ),
       .io_input( T25 ),
       .io_output( CircularPeekQueue_io_output )
  );
  CircularPeekQueue_1 CircularPeekQueue_1(.clk(clk), .reset(reset),
       .io_writeEnable( T23 ),
       .io_nextBlock( T21 ),
       .io_input( T16 ),
       .io_output( CircularPeekQueue_1_io_output )
  );
  CircularPeekQueue_1 CircularPeekQueue_2(.clk(clk), .reset(reset),
       .io_writeEnable( T12 ),
       .io_nextBlock( T9 ),
       .io_input( T4 ),
       .io_output( CircularPeekQueue_2_io_output )
  );
  WrappingCounter_0 inputSelectCounter(
       .io_enable( R3 ),
       .io_value( inputSelectCounter_io_value )
  );
  WrappingCounter_1 inputSelectCounter_1(
       .io_enable( R2 ),
       .io_value( inputSelectCounter_1_io_value )
  );
  WrappingCounter_2 inputSelectCounter_2(
       .io_enable( R1 ),
       .io_value( inputSelectCounter_2_io_value )
  );
  WrappingCounter_0 queueOutputSelectCounters(
       .io_enable( signalNewPeekBlock ),
       .io_value( queueOutputSelectCounters_io_value )
  );
  WrappingCounter_1 queueOutputSelectCounters_1(
       .io_enable( signalNewPeekBlock ),
       .io_value( queueOutputSelectCounters_1_io_value )
  );
  WrappingCounter_2 queueOutputSelectCounters_2(
       .io_enable( signalNewPeekBlock ),
       .io_value( queueOutputSelectCounters_2_io_value )
  );
  WrappingCounter_0 outputSelectCounters(
       .io_enable( signalNewPeekBlock ),
       .io_value( outputSelectCounters_io_value )
  );
  WrappingCounter_1 outputSelectCounters_1(
       .io_enable( signalNewPeekBlock ),
       .io_value( outputSelectCounters_1_io_value )
  );
  WrappingCounter_2 outputSelectCounters_2(
       .io_enable( signalNewPeekBlock ),
       .io_value( outputSelectCounters_2_io_value )
  );

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else begin
      R1 <= io_prevDone;
    end
    if(reset) begin
      R2 <= 1'h0;
    end else begin
      R2 <= io_prevDone;
    end
    if(reset) begin
      R3 <= 1'h0;
    end else begin
      R3 <= io_prevDone;
    end
    if(reset) begin
      signalBitBuffersFull <= 1'h0;
    end else begin
      signalBitBuffersFull <= T15;
    end
    if(reset) begin
      R34 <= 1'h0;
    end else begin
      R34 <= io_prevDone;
    end
    if(reset) begin
      R35 <= 1'h0;
    end else begin
      R35 <= io_prevDone;
    end
    if(reset) begin
      R51 <= 1'h0;
    end else begin
      R51 <= signalNewPeekBlock;
    end
  end
endmodule

module UpDownCounter_3(input clk, input reset,
    input  io_up,
    input  io_down,
    output[3:0] io_value
);

  reg [3:0] reg_;
  wire[3:0] T10;
  wire[3:0] T0;
  wire[3:0] T1;
  wire[3:0] T2;
  wire T3;
  wire T4;
  wire T5;
  wire[3:0] T6;
  wire T7;
  wire T8;
  wire T9;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    reg_ = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = reg_;
  assign T10 = reset ? 4'h0 : T0;
  assign T0 = T7 ? T6 : T1;
  assign T1 = T3 ? T2 : reg_;
  assign T2 = reg_ + 4'h3;
  assign T3 = T4 & io_up;
  assign T4 = T5 ^ 1'h1;
  assign T5 = io_up & io_down;
  assign T6 = reg_ - 4'h1;
  assign T7 = T8 & io_down;
  assign T8 = T9 ^ 1'h1;
  assign T9 = T5 | io_up;

  always @(posedge clk) begin
    if(reset) begin
      reg_ <= 4'h0;
    end else if(T7) begin
      reg_ <= T6;
    end else if(T3) begin
      reg_ <= T2;
    end
  end
endmodule

module WrappingCounter_11(input clk, input reset,
    input  io_enable,
    output[2:0] io_value
);

  reg [2:0] R0;
  wire[2:0] T11;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire T5;
  wire T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire T9;
  wire T10;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = R0;
  assign T11 = reset ? 3'h2 : T1;
  assign T1 = T9 ? T8 : T2;
  assign T2 = T5 ? T3 : R0;
  assign T3 = T4 - 3'h3;
  assign T4 = R0 + 3'h1;
  assign T5 = io_enable & T6;
  assign T6 = 3'h3 <= T7;
  assign T7 = R0 + 3'h1;
  assign T8 = R0 + 3'h1;
  assign T9 = io_enable & T10;
  assign T10 = T6 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R0 <= 3'h2;
    end else if(T9) begin
      R0 <= T8;
    end else if(T5) begin
      R0 <= T3;
    end
  end
endmodule

module WrappingCounter_12(input clk, input reset,
    input  io_enable,
    output[2:0] io_value
);

  reg [2:0] R0;
  wire[2:0] T11;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire T5;
  wire T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire T9;
  wire T10;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = R0;
  assign T11 = reset ? 3'h0 : T1;
  assign T1 = T9 ? T8 : T2;
  assign T2 = T5 ? T3 : R0;
  assign T3 = T4 - 3'h3;
  assign T4 = R0 + 3'h2;
  assign T5 = io_enable & T6;
  assign T6 = 3'h3 <= T7;
  assign T7 = R0 + 3'h2;
  assign T8 = R0 + 3'h2;
  assign T9 = io_enable & T10;
  assign T10 = T6 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R0 <= 3'h0;
    end else if(T9) begin
      R0 <= T8;
    end else if(T5) begin
      R0 <= T3;
    end
  end
endmodule

module WrappingCounter_13(input clk, input reset,
    input  io_enable,
    output[2:0] io_value
);

  reg [2:0] R0;
  wire[2:0] T11;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire T5;
  wire T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire T9;
  wire T10;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = R0;
  assign T11 = reset ? 3'h1 : T1;
  assign T1 = T9 ? T8 : T2;
  assign T2 = T5 ? T3 : R0;
  assign T3 = T4 - 3'h3;
  assign T4 = R0 + 3'h2;
  assign T5 = io_enable & T6;
  assign T6 = 3'h3 <= T7;
  assign T7 = R0 + 3'h2;
  assign T8 = R0 + 3'h2;
  assign T9 = io_enable & T10;
  assign T10 = T6 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R0 <= 3'h1;
    end else if(T9) begin
      R0 <= T8;
    end else if(T5) begin
      R0 <= T3;
    end
  end
endmodule

module WrappingCounter_14(input clk, input reset,
    input  io_enable,
    output[2:0] io_value
);

  reg [2:0] R0;
  wire[2:0] T11;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire T5;
  wire T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire T9;
  wire T10;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_value = R0;
  assign T11 = reset ? 3'h2 : T1;
  assign T1 = T9 ? T8 : T2;
  assign T2 = T5 ? T3 : R0;
  assign T3 = T4 - 3'h3;
  assign T4 = R0 + 3'h2;
  assign T5 = io_enable & T6;
  assign T6 = 3'h3 <= T7;
  assign T7 = R0 + 3'h2;
  assign T8 = R0 + 3'h2;
  assign T9 = io_enable & T10;
  assign T10 = T6 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R0 <= 3'h2;
    end else if(T9) begin
      R0 <= T8;
    end else if(T5) begin
      R0 <= T3;
    end
  end
endmodule

module GearBox_2(input clk, input reset,
    input  io_xsIn_2,
    input  io_xsIn_1,
    input  io_xsIn_0,
    input  io_validIn,
    input  io_prevDone,
    input  io_prevStart,
    output io_ready,
    input  io_nextReady,
    output io_startNext,
    output[15:0] io_xsOut_0
);

  wire signalNewPeekBlock;
  wire T0;
  reg  R1;
  wire T42;
  reg  R2;
  wire T43;
  reg  R3;
  wire T44;
  wire[15:0] T4;
  wire[15:0] T5;
  wire T6;
  wire[1:0] T7;
  wire T8;
  wire T9;
  reg  T10;
  wire[1:0] T45;
  wire T12;
  reg  T13;
  reg  signalBitBuffersFull;
  wire T46;
  wire T15;
  wire signalResetBitBuffers;
  wire[15:0] T16;
  wire[15:0] T17;
  wire T18;
  wire[1:0] T19;
  wire[1:0] T47;
  wire T20;
  wire T21;
  reg  T22;
  wire[1:0] T48;
  wire T23;
  reg  T24;
  wire[1:0] T49;
  wire[15:0] T25;
  wire[15:0] T26;
  wire T27;
  wire[1:0] T28;
  wire[1:0] T50;
  wire T29;
  wire T30;
  reg  T31;
  wire[1:0] T51;
  wire T32;
  reg  T33;
  wire[1:0] T52;
  reg  R34;
  wire T53;
  reg  R35;
  wire T54;
  wire[15:0] T36;
  wire[15:0] T37;
  wire T38;
  wire[1:0] T39;
  wire[1:0] T55;
  wire T40;
  reg  R41;
  wire T56;
  wire hasEnoughEmptyBlocks;
  wire[3:0] reservedBlocks;
  wire[3:0] T57;
  wire[15:0] BitToWord_io_word;
  wire[15:0] BitToWord_1_io_word;
  wire[15:0] BitToWord_2_io_word;
  wire[2:0] fillingBlock_io_value;
  wire[3:0] bitCounter_io_value;
  wire[3:0] blocksReady_io_value;
  wire inputSelectCounter_io_value;
  wire inputSelectCounter_1_io_value;
  wire[1:0] inputSelectCounter_2_io_value;
  wire[2:0] queueOutputSelectCounters_io_value;
  wire[2:0] outputSelectCounters_io_value;
  wire[2:0] outputSelectCounters_1_io_value;
  wire[2:0] outputSelectCounters_2_io_value;
  wire[15:0] CircularPeekQueue_io_output;
  wire[15:0] CircularPeekQueue_1_io_output;
  wire[15:0] CircularPeekQueue_2_io_output;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R2 = {1{$random}};
    R3 = {1{$random}};
    signalBitBuffersFull = {1{$random}};
    R34 = {1{$random}};
    R35 = {1{$random}};
    R41 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign signalNewPeekBlock = io_nextReady & T0;
  assign T0 = 4'h1 <= blocksReady_io_value;
  assign T42 = reset ? 1'h0 : io_prevDone;
  assign T43 = reset ? 1'h0 : io_prevDone;
  assign T44 = reset ? 1'h0 : io_prevDone;
  assign T4 = T8 ? BitToWord_2_io_word : T5;
  assign T5 = T6 ? BitToWord_1_io_word : BitToWord_io_word;
  assign T6 = T7[0];
  assign T7 = inputSelectCounter_2_io_value;
  assign T8 = T7[1];
  assign T9 = signalNewPeekBlock & T10;
  always @(*) case (T45)
    0: T10 = 1'h1;
    1: T10 = 1'h0;
    2: T10 = 1'h0;
    default: begin
      T10 = 1'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T10 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T45 = outputSelectCounters_2_io_value[1:0];
  assign T12 = signalBitBuffersFull & T13;
  always @(*) case (inputSelectCounter_2_io_value)
    0: T13 = 1'h1;
    1: T13 = 1'h1;
    2: T13 = 1'h1;
    default: begin
      T13 = 1'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T13 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T46 = reset ? 1'h0 : T15;
  assign T15 = io_validIn & signalResetBitBuffers;
  assign signalResetBitBuffers = bitCounter_io_value == 4'hf;
  assign T16 = T20 ? BitToWord_2_io_word : T17;
  assign T17 = T18 ? BitToWord_1_io_word : BitToWord_io_word;
  assign T18 = T19[0];
  assign T19 = T47;
  assign T47 = {1'h0, inputSelectCounter_1_io_value};
  assign T20 = T19[1];
  assign T21 = signalNewPeekBlock & T22;
  always @(*) case (T48)
    0: T22 = 1'h1;
    1: T22 = 1'h0;
    2: T22 = 1'h0;
    default: begin
      T22 = 1'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T22 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T48 = outputSelectCounters_1_io_value[1:0];
  assign T23 = signalBitBuffersFull & T24;
  always @(*) case (T49)
    0: T24 = 1'h1;
    1: T24 = 1'h1;
    2: T24 = 1'h1;
    default: begin
      T24 = 1'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T24 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T49 = {1'h0, inputSelectCounter_1_io_value};
  assign T25 = T29 ? BitToWord_2_io_word : T26;
  assign T26 = T27 ? BitToWord_1_io_word : BitToWord_io_word;
  assign T27 = T28[0];
  assign T28 = T50;
  assign T50 = {1'h0, inputSelectCounter_io_value};
  assign T29 = T28[1];
  assign T30 = signalNewPeekBlock & T31;
  always @(*) case (T51)
    0: T31 = 1'h1;
    1: T31 = 1'h0;
    2: T31 = 1'h0;
    default: begin
      T31 = 1'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T31 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T51 = outputSelectCounters_io_value[1:0];
  assign T32 = signalBitBuffersFull & T33;
  always @(*) case (T52)
    0: T33 = 1'h1;
    1: T33 = 1'h1;
    2: T33 = 1'h1;
    default: begin
      T33 = 1'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T33 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T52 = {1'h0, inputSelectCounter_io_value};
  assign T53 = reset ? 1'h0 : io_prevDone;
  assign T54 = reset ? 1'h0 : io_prevDone;
  assign io_xsOut_0 = T36;
  assign T36 = T40 ? CircularPeekQueue_2_io_output : T37;
  assign T37 = T38 ? CircularPeekQueue_1_io_output : CircularPeekQueue_io_output;
  assign T38 = T39[0];
  assign T39 = T55;
  assign T55 = queueOutputSelectCounters_io_value[1:0];
  assign T40 = T39[1];
  assign io_startNext = R41;
  assign T56 = reset ? 1'h0 : signalNewPeekBlock;
  assign io_ready = hasEnoughEmptyBlocks;
  assign hasEnoughEmptyBlocks = reservedBlocks <= 4'h5;
  assign reservedBlocks = blocksReady_io_value + T57;
  assign T57 = {1'h0, fillingBlock_io_value};
  BitToWord_1 BitToWord(.clk(clk),
       .io_enable( io_validIn ),
       .io_bit( io_xsIn_0 ),
       .io_word( BitToWord_io_word )
  );
  BitToWord_1 BitToWord_1(.clk(clk),
       .io_enable( io_validIn ),
       .io_bit( io_xsIn_1 ),
       .io_word( BitToWord_1_io_word )
  );
  BitToWord_1 BitToWord_2(.clk(clk),
       .io_enable( io_validIn ),
       .io_bit( io_xsIn_2 ),
       .io_word( BitToWord_2_io_word )
  );
  AsyncUpDownCounter_1 fillingBlock(.clk(clk), .reset(reset),
       .io_up( io_prevStart ),
       .io_down( R35 ),
       .io_value( fillingBlock_io_value )
  );
  Counter_2 bitCounter(.clk(clk), .reset(reset),
       .io_enable( io_validIn ),
       .io_rst( signalResetBitBuffers ),
       .io_value( bitCounter_io_value )
  );
  UpDownCounter_3 blocksReady(.clk(clk), .reset(reset),
       .io_up( R34 ),
       .io_down( signalNewPeekBlock ),
       .io_value( blocksReady_io_value )
  );
  CircularPeekQueue_1 CircularPeekQueue(.clk(clk), .reset(reset),
       .io_writeEnable( T32 ),
       .io_nextBlock( T30 ),
       .io_input( T25 ),
       .io_output( CircularPeekQueue_io_output )
  );
  CircularPeekQueue_1 CircularPeekQueue_1(.clk(clk), .reset(reset),
       .io_writeEnable( T23 ),
       .io_nextBlock( T21 ),
       .io_input( T16 ),
       .io_output( CircularPeekQueue_1_io_output )
  );
  CircularPeekQueue_1 CircularPeekQueue_2(.clk(clk), .reset(reset),
       .io_writeEnable( T12 ),
       .io_nextBlock( T9 ),
       .io_input( T4 ),
       .io_output( CircularPeekQueue_2_io_output )
  );
  WrappingCounter_0 inputSelectCounter(
       .io_enable( R3 ),
       .io_value( inputSelectCounter_io_value )
  );
  WrappingCounter_1 inputSelectCounter_1(
       .io_enable( R2 ),
       .io_value( inputSelectCounter_1_io_value )
  );
  WrappingCounter_2 inputSelectCounter_2(
       .io_enable( R1 ),
       .io_value( inputSelectCounter_2_io_value )
  );
  WrappingCounter_11 queueOutputSelectCounters(.clk(clk), .reset(reset),
       .io_enable( signalNewPeekBlock ),
       .io_value( queueOutputSelectCounters_io_value )
  );
  WrappingCounter_12 outputSelectCounters(.clk(clk), .reset(reset),
       .io_enable( signalNewPeekBlock ),
       .io_value( outputSelectCounters_io_value )
  );
  WrappingCounter_13 outputSelectCounters_1(.clk(clk), .reset(reset),
       .io_enable( signalNewPeekBlock ),
       .io_value( outputSelectCounters_1_io_value )
  );
  WrappingCounter_14 outputSelectCounters_2(.clk(clk), .reset(reset),
       .io_enable( signalNewPeekBlock ),
       .io_value( outputSelectCounters_2_io_value )
  );

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else begin
      R1 <= io_prevDone;
    end
    if(reset) begin
      R2 <= 1'h0;
    end else begin
      R2 <= io_prevDone;
    end
    if(reset) begin
      R3 <= 1'h0;
    end else begin
      R3 <= io_prevDone;
    end
    if(reset) begin
      signalBitBuffersFull <= 1'h0;
    end else begin
      signalBitBuffersFull <= T15;
    end
    if(reset) begin
      R34 <= 1'h0;
    end else begin
      R34 <= io_prevDone;
    end
    if(reset) begin
      R35 <= 1'h0;
    end else begin
      R35 <= io_prevDone;
    end
    if(reset) begin
      R41 <= 1'h0;
    end else begin
      R41 <= signalNewPeekBlock;
    end
  end
endmodule

module Net(input clk, input reset,
    output io_ready,
    input  io_start,
    input [15:0] io_xsIn_3,
    input [15:0] io_xsIn_2,
    input [15:0] io_xsIn_1,
    input [15:0] io_xsIn_0,
    output io_xsOut_0,
    output io_xsOutValid,
    output io_done,
    input  io_pipeReady
);

  wire Warp_io_ready;
  wire Warp_io_startOut;
  wire Warp_io_xOut_3;
  wire Warp_io_xOut_2;
  wire Warp_io_xOut_1;
  wire Warp_io_xOut_0;
  wire Warp_io_xOutValid;
  wire Warp_io_done;
  wire Warp_1_io_ready;
  wire Warp_1_io_startOut;
  wire Warp_1_io_xOut_2;
  wire Warp_1_io_xOut_1;
  wire Warp_1_io_xOut_0;
  wire Warp_1_io_xOutValid;
  wire Warp_1_io_done;
  wire Warp_2_io_ready;
  wire Warp_2_io_startOut;
  wire Warp_2_io_xOut_2;
  wire Warp_2_io_xOut_1;
  wire Warp_2_io_xOut_0;
  wire Warp_2_io_xOutValid;
  wire Warp_2_io_done;
  wire Warp_3_io_ready;
  wire Warp_3_io_xOut_0;
  wire Warp_3_io_xOutValid;
  wire Warp_3_io_done;
  wire GearBox_io_ready;
  wire GearBox_io_startNext;
  wire[15:0] GearBox_io_xsOut_2;
  wire[15:0] GearBox_io_xsOut_1;
  wire[15:0] GearBox_io_xsOut_0;
  wire GearBox_1_io_ready;
  wire GearBox_1_io_startNext;
  wire[15:0] GearBox_1_io_xsOut_2;
  wire[15:0] GearBox_1_io_xsOut_1;
  wire[15:0] GearBox_1_io_xsOut_0;
  wire GearBox_2_io_ready;
  wire GearBox_2_io_startNext;
  wire[15:0] GearBox_2_io_xsOut_0;


  assign io_done = Warp_3_io_done;
  assign io_xsOutValid = Warp_3_io_xOutValid;
  assign io_xsOut_0 = Warp_3_io_xOut_0;
  assign io_ready = Warp_io_ready;
  Warp_0 Warp(.clk(clk), .reset(reset),
       .io_xIn_3( io_xsIn_3 ),
       .io_xIn_2( io_xsIn_2 ),
       .io_xIn_1( io_xsIn_1 ),
       .io_xIn_0( io_xsIn_0 ),
       .io_start( io_start ),
       .io_ready( Warp_io_ready ),
       .io_startOut( Warp_io_startOut ),
       .io_xOut_3( Warp_io_xOut_3 ),
       .io_xOut_2( Warp_io_xOut_2 ),
       .io_xOut_1( Warp_io_xOut_1 ),
       .io_xOut_0( Warp_io_xOut_0 ),
       .io_xOutValid( Warp_io_xOutValid ),
       .io_pipeReady( GearBox_io_ready ),
       .io_done( Warp_io_done )
  );
  Warp_1 Warp_1(.clk(clk), .reset(reset),
       .io_xIn_2( GearBox_io_xsOut_2 ),
       .io_xIn_1( GearBox_io_xsOut_1 ),
       .io_xIn_0( GearBox_io_xsOut_0 ),
       .io_start( GearBox_io_startNext ),
       .io_ready( Warp_1_io_ready ),
       .io_startOut( Warp_1_io_startOut ),
       .io_xOut_2( Warp_1_io_xOut_2 ),
       .io_xOut_1( Warp_1_io_xOut_1 ),
       .io_xOut_0( Warp_1_io_xOut_0 ),
       .io_xOutValid( Warp_1_io_xOutValid ),
       .io_pipeReady( GearBox_1_io_ready ),
       .io_done( Warp_1_io_done )
  );
  Warp_2 Warp_2(.clk(clk), .reset(reset),
       .io_xIn_2( GearBox_1_io_xsOut_2 ),
       .io_xIn_1( GearBox_1_io_xsOut_1 ),
       .io_xIn_0( GearBox_1_io_xsOut_0 ),
       .io_start( GearBox_1_io_startNext ),
       .io_ready( Warp_2_io_ready ),
       .io_startOut( Warp_2_io_startOut ),
       .io_xOut_2( Warp_2_io_xOut_2 ),
       .io_xOut_1( Warp_2_io_xOut_1 ),
       .io_xOut_0( Warp_2_io_xOut_0 ),
       .io_xOutValid( Warp_2_io_xOutValid ),
       .io_pipeReady( GearBox_2_io_ready ),
       .io_done( Warp_2_io_done )
  );
  Warp_3 Warp_3(.clk(clk), .reset(reset),
       .io_xIn_0( GearBox_2_io_xsOut_0 ),
       .io_start( GearBox_2_io_startNext ),
       .io_ready( Warp_3_io_ready ),
       //.io_startOut(  )
       .io_xOut_0( Warp_3_io_xOut_0 ),
       .io_xOutValid( Warp_3_io_xOutValid ),
       .io_pipeReady( io_pipeReady ),
       .io_done( Warp_3_io_done )
  );
  GearBox_0 GearBox(.clk(clk), .reset(reset),
       .io_xsIn_3( Warp_io_xOut_3 ),
       .io_xsIn_2( Warp_io_xOut_2 ),
       .io_xsIn_1( Warp_io_xOut_1 ),
       .io_xsIn_0( Warp_io_xOut_0 ),
       .io_validIn( Warp_io_xOutValid ),
       .io_prevDone( Warp_io_done ),
       .io_prevStart( Warp_io_startOut ),
       .io_ready( GearBox_io_ready ),
       .io_nextReady( Warp_1_io_ready ),
       .io_startNext( GearBox_io_startNext ),
       .io_xsOut_2( GearBox_io_xsOut_2 ),
       .io_xsOut_1( GearBox_io_xsOut_1 ),
       .io_xsOut_0( GearBox_io_xsOut_0 )
  );
  GearBox_1 GearBox_1(.clk(clk), .reset(reset),
       .io_xsIn_2( Warp_1_io_xOut_2 ),
       .io_xsIn_1( Warp_1_io_xOut_1 ),
       .io_xsIn_0( Warp_1_io_xOut_0 ),
       .io_validIn( Warp_1_io_xOutValid ),
       .io_prevDone( Warp_1_io_done ),
       .io_prevStart( Warp_1_io_startOut ),
       .io_ready( GearBox_1_io_ready ),
       .io_nextReady( Warp_2_io_ready ),
       .io_startNext( GearBox_1_io_startNext ),
       .io_xsOut_2( GearBox_1_io_xsOut_2 ),
       .io_xsOut_1( GearBox_1_io_xsOut_1 ),
       .io_xsOut_0( GearBox_1_io_xsOut_0 )
  );
  GearBox_2 GearBox_2(.clk(clk), .reset(reset),
       .io_xsIn_2( Warp_2_io_xOut_2 ),
       .io_xsIn_1( Warp_2_io_xOut_1 ),
       .io_xsIn_0( Warp_2_io_xOut_0 ),
       .io_validIn( Warp_2_io_xOutValid ),
       .io_prevDone( Warp_2_io_done ),
       .io_prevStart( Warp_2_io_startOut ),
       .io_ready( GearBox_2_io_ready ),
       .io_nextReady( Warp_3_io_ready ),
       .io_startNext( GearBox_2_io_startNext ),
       .io_xsOut_0( GearBox_2_io_xsOut_0 )
  );
endmodule

module BitToWord_0(input clk,
    input  io_enable,
    input  io_bit,
    output[9:0] io_word
);

  wire[9:0] T0;
  reg  R1;
  wire T2;
  reg  R3;
  wire T4;
  reg  R5;
  wire T6;
  reg  R7;
  wire T8;
  reg  R9;
  wire T10;
  reg  R11;
  wire T12;
  reg  R13;
  wire T14;
  reg  R15;
  wire T16;
  reg  R17;
  wire T18;
  reg  R19;
  wire T20;
  wire[8:0] T21;
  wire[7:0] T22;
  wire[6:0] T23;
  wire[5:0] T24;
  wire[4:0] T25;
  wire[3:0] T26;
  wire[2:0] T27;
  wire[1:0] T28;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R3 = {1{$random}};
    R5 = {1{$random}};
    R7 = {1{$random}};
    R9 = {1{$random}};
    R11 = {1{$random}};
    R13 = {1{$random}};
    R15 = {1{$random}};
    R17 = {1{$random}};
    R19 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_word = T0;
  assign T0 = {T21, R1};
  assign T2 = io_enable ? R3 : R1;
  assign T4 = io_enable ? R5 : R3;
  assign T6 = io_enable ? R7 : R5;
  assign T8 = io_enable ? R9 : R7;
  assign T10 = io_enable ? R11 : R9;
  assign T12 = io_enable ? R13 : R11;
  assign T14 = io_enable ? R15 : R13;
  assign T16 = io_enable ? R17 : R15;
  assign T18 = io_enable ? R19 : R17;
  assign T20 = io_enable ? io_bit : R19;
  assign T21 = {T22, R3};
  assign T22 = {T23, R5};
  assign T23 = {T24, R7};
  assign T24 = {T25, R9};
  assign T25 = {T26, R11};
  assign T26 = {T27, R13};
  assign T27 = {T28, R15};
  assign T28 = {R19, R17};

  always @(posedge clk) begin
    if(io_enable) begin
      R1 <= R3;
    end
    if(io_enable) begin
      R3 <= R5;
    end
    if(io_enable) begin
      R5 <= R7;
    end
    if(io_enable) begin
      R7 <= R9;
    end
    if(io_enable) begin
      R9 <= R11;
    end
    if(io_enable) begin
      R11 <= R13;
    end
    if(io_enable) begin
      R13 <= R15;
    end
    if(io_enable) begin
      R15 <= R17;
    end
    if(io_enable) begin
      R17 <= R19;
    end
    if(io_enable) begin
      R19 <= io_bit;
    end
  end
endmodule

module Deinterleaver(input clk, input reset,
    output io_oneBitPerCore_ready,
    input  io_oneBitPerCore_valid,
    input  io_oneBitPerCore_bits,
    input  io_oneHotOut_ready,
    output io_oneHotOut_valid,
    output[9:0] io_oneHotOut_bits,
    input  io_doneIn
);

  reg [9:0] regsBuf_0;
  wire[9:0] T7;
  wire[9:0] T0;
  reg  doneDelay;
  wire T8;
  reg  send;
  wire T9;
  wire T1;
  wire T2;
  wire T3;
  reg  count;
  wire T10;
  wire T4;
  wire T5;
  wire T6;
  wire[9:0] BitToWord_io_word;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    regsBuf_0 = {1{$random}};
    doneDelay = {1{$random}};
    send = {1{$random}};
    count = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_oneHotOut_bits = regsBuf_0;
  assign T7 = reset ? 10'h0 : T0;
  assign T0 = doneDelay ? BitToWord_io_word : regsBuf_0;
  assign T8 = reset ? 1'h0 : io_doneIn;
  assign io_oneHotOut_valid = send;
  assign T9 = reset ? 1'h0 : T1;
  assign T1 = T2 ? doneDelay : send;
  assign T2 = doneDelay | T3;
  assign T3 = count == 1'h0;
  assign T10 = reset ? 1'h0 : T4;
  assign T4 = T5 ? 1'h0 : count;
  assign T5 = send & T6;
  assign T6 = count == 1'h0;
  assign io_oneBitPerCore_ready = io_oneHotOut_ready;
  BitToWord_0 BitToWord(.clk(clk),
       .io_enable( io_oneBitPerCore_valid ),
       .io_bit( io_oneBitPerCore_bits ),
       .io_word( BitToWord_io_word )
  );

  always @(posedge clk) begin
    if(reset) begin
      regsBuf_0 <= 10'h0;
    end else if(doneDelay) begin
      regsBuf_0 <= BitToWord_io_word;
    end
    if(reset) begin
      doneDelay <= 1'h0;
    end else begin
      doneDelay <= io_doneIn;
    end
    if(reset) begin
      send <= 1'h0;
    end else if(T2) begin
      send <= doneDelay;
    end
    if(reset) begin
      count <= 1'h0;
    end else if(T5) begin
      count <= 1'h0;
    end
  end
endmodule

module Pacman(input clk, input reset,
    output io_inDataStream_ready,
    input  io_inDataStream_valid,
    input [7:0] io_inDataStream_bits,
    input  io_digitOut_ready,
    output io_digitOut_valid,
    output[3:0] io_digitOut_bits
);

  wire[3:0] T1;
  wire[2:0] T2;
  wire[1:0] T3;
  wire T4;
  wire[1:0] T5;
  wire[1:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[7:0] T9;
  wire[7:0] T10;
  wire[1:0] T11;
  wire[3:0] T12;
  wire[1:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire widthConverter_io_wordIn_ready;
  wire widthConverter_io_wordOut_valid;
  wire[15:0] widthConverter_io_wordOut_bits;
  wire deinterleaver_io_oneBitPerCore_ready;
  wire deinterleaver_io_oneHotOut_valid;
  wire[9:0] deinterleaver_io_oneHotOut_bits;
  wire interleaver_io_wordIn_ready;
  wire[15:0] interleaver_io_interleavedOut_3;
  wire[15:0] interleaver_io_interleavedOut_2;
  wire[15:0] interleaver_io_interleavedOut_1;
  wire[15:0] interleaver_io_interleavedOut_0;
  wire interleaver_io_startOut;
  wire net_io_ready;
  wire net_io_xsOut_0;
  wire net_io_xsOutValid;
  wire net_io_done;


  assign io_digitOut_bits = T1;
  assign T1 = {T16, T2};
  assign T2 = {T15, T3};
  assign T3 = {T14, T4};
  assign T4 = T5[1];
  assign T5 = T13 | T6;
  assign T6 = T7[1:0];
  assign T7 = T12 | T8;
  assign T8 = T9[3:0];
  assign T9 = T11 | T10;
  assign T10 = deinterleaver_io_oneHotOut_bits[7:0];
  assign T11 = deinterleaver_io_oneHotOut_bits[9:8];
  assign T12 = T9[7:4];
  assign T13 = T7[3:2];
  assign T14 = T13 != 2'h0;
  assign T15 = T12 != 4'h0;
  assign T16 = T11 != 2'h0;
  assign io_digitOut_valid = deinterleaver_io_oneHotOut_valid;
  assign io_inDataStream_ready = widthConverter_io_wordIn_ready;
  WidthConverter widthConverter(.clk(clk), .reset(reset),
       .io_wordIn_ready( widthConverter_io_wordIn_ready ),
       .io_wordIn_valid( io_inDataStream_valid ),
       .io_wordIn_bits( io_inDataStream_bits ),
       .io_wordOut_ready( interleaver_io_wordIn_ready ),
       .io_wordOut_valid( widthConverter_io_wordOut_valid ),
       .io_wordOut_bits( widthConverter_io_wordOut_bits )
  );
  Interleaver interleaver(.clk(clk), .reset(reset),
       .io_wordIn_ready( interleaver_io_wordIn_ready ),
       .io_wordIn_valid( widthConverter_io_wordOut_valid ),
       .io_wordIn_bits( widthConverter_io_wordOut_bits ),
       .io_interleavedOut_3( interleaver_io_interleavedOut_3 ),
       .io_interleavedOut_2( interleaver_io_interleavedOut_2 ),
       .io_interleavedOut_1( interleaver_io_interleavedOut_1 ),
       .io_interleavedOut_0( interleaver_io_interleavedOut_0 ),
       .io_startOut( interleaver_io_startOut ),
       .io_pipeReady( net_io_ready )
  );
  Net net(.clk(clk), .reset(reset),
       .io_ready( net_io_ready ),
       .io_start( interleaver_io_startOut ),
       .io_xsIn_3( interleaver_io_interleavedOut_3 ),
       .io_xsIn_2( interleaver_io_interleavedOut_2 ),
       .io_xsIn_1( interleaver_io_interleavedOut_1 ),
       .io_xsIn_0( interleaver_io_interleavedOut_0 ),
       .io_xsOut_0( net_io_xsOut_0 ),
       .io_xsOutValid( net_io_xsOutValid ),
       .io_done( net_io_done ),
       .io_pipeReady( deinterleaver_io_oneBitPerCore_ready )
  );
  Deinterleaver deinterleaver(.clk(clk), .reset(reset),
       .io_oneBitPerCore_ready( deinterleaver_io_oneBitPerCore_ready ),
       .io_oneBitPerCore_valid( net_io_xsOutValid ),
       .io_oneBitPerCore_bits( net_io_xsOut_0 ),
       .io_oneHotOut_ready( io_digitOut_ready ),
       .io_oneHotOut_valid( deinterleaver_io_oneHotOut_valid ),
       .io_oneHotOut_bits( deinterleaver_io_oneHotOut_bits ),
       .io_doneIn( net_io_done )
  );
endmodule

module PacmanWrapper(input ulpi_clk, input clk, input reset,
    output io_usb_data_ready,
    input  io_usb_data_valid,
    input [7:0] io_usb_data_bits,
    input  io_net_result_ready,
    output io_net_result_valid,
    output[3:0] io_net_result_bits
);

  wire AsyncFifo_inst_io_enq_ready;
  wire AsyncFifo_inst_io_deq_valid;
  wire[7:0] AsyncFifo_inst_io_deq_bits;
  wire Pacman_inst_io_inDataStream_ready;
  wire Pacman_inst_io_digitOut_valid;
  wire[3:0] Pacman_inst_io_digitOut_bits;


  assign io_net_result_bits = Pacman_inst_io_digitOut_bits;
  assign io_net_result_valid = Pacman_inst_io_digitOut_valid;
  assign io_usb_data_ready = AsyncFifo_inst_io_enq_ready;
  AsyncFifo AsyncFifo_inst(.ulpi_clk(ulpi_clk), .clk(clk), .reset(reset),
       .io_enq_ready( AsyncFifo_inst_io_enq_ready ),
       .io_enq_valid( io_usb_data_valid ),
       .io_enq_bits( io_usb_data_bits ),
       .io_deq_ready( Pacman_inst_io_inDataStream_ready ),
       .io_deq_valid( AsyncFifo_inst_io_deq_valid ),
       .io_deq_bits( AsyncFifo_inst_io_deq_bits )
       //.io_count(  )
  );
  Pacman Pacman_inst(.clk(clk), .reset(reset),
       .io_inDataStream_ready( Pacman_inst_io_inDataStream_ready ),
       .io_inDataStream_valid( AsyncFifo_inst_io_deq_valid ),
       .io_inDataStream_bits( AsyncFifo_inst_io_deq_bits ),
       .io_digitOut_ready( io_net_result_ready ),
       .io_digitOut_valid( Pacman_inst_io_digitOut_valid ),
       .io_digitOut_bits( Pacman_inst_io_digitOut_bits )
  );
endmodule

